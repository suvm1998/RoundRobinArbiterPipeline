module arbiter(a, b, c, d, clk, rst, out);
wire [1:0] _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
input a;
input b;
input c;
input clk;
wire [1:0] counter;
input d;
output out;
input rst;
NOT _16_ (.A(b),.Y(_03_));
NOR _21_ (.A(_05_),.B(_07_),.Y(_08_));
NAND _25_ (.A(_00_[0]),.B(_11_),.Y(_12_));
NAND _26_ (.A(_08_),.B(_12_),.Y(_01_));
DFF _29_ (.C(clk),.D(_00_[0]),.Q(counter[0]));
DFF _30_ (.C(clk),.D(_00_[1]),.Q(counter[1]));
DFF _31_ (.C(clk),.D(_01_),.Q(out));
input _0_0_;
NOT _14_ (.A(counter[0]),.Y(_0_0_));
DFF _0_0_0_ (.C(clk),.D(_0_0_),.Y(_00_[0]));
input _1_1_;
NOR _20_ (.A(_00_[0]),.B(_06_),.Y(_1_1_));
DFF _1_1_1_ (.C(clk),.D(_1_1_),.Y(_07_));
input _2_2_;
NAND _27_ (.A(_00_[0]),.B(counter[1]),.Y(_2_2_));
DFF _2_2_2_ (.C(clk),.D(_2_2_),.Y(_13_));
input _3_3_;
NOR _23_ (.A(counter[1]),.B(a),.Y(_3_3_));
DFF _3_3_3_ (.C(clk),.D(_3_3_),.Y(_10_));
input _4_4_;
NOR _22_ (.A(_02_),.B(c),.Y(_4_4_));
DFF _4_4_4_ (.C(clk),.D(_4_4_),.Y(_09_));
input _5_5_;
NAND _17_ (.A(counter[0]),.B(_02_),.Y(_5_5_));
DFF _5_5_5_ (.C(clk),.D(_5_5_),.Y(_04_));
input _6_6_;
NAND _19_ (.A(counter[1]),.B(d),.Y(_6_6_));
DFF _6_6_6_ (.C(clk),.D(_6_6_),.Y(_06_));
input _7_7_;
NOT _15_ (.A(counter[1]),.Y(_7_7_));
DFF _7_7_7_ (.C(clk),.D(_7_7_),.Y(_02_));
input _8_8_;
NOR _24_ (.A(_09_),.B(_10_),.Y(_8_8_));
DFF _8_8_8_ (.C(clk),.D(_8_8_),.Y(_11_));
input _9_9_;
NAND _28_ (.A(_04_),.B(_13_),.Y(_9_9_));
DFF _9_9_9_ (.C(clk),.D(_9_9_),.Y(_00_[1]));
input _10_10_;
NOR _18_ (.A(_03_),.B(_04_),.Y(_10_10_));
DFF _10_10_10_ (.C(clk),.D(_10_10_),.Y(_05_));

endmodule

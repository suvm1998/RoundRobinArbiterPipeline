module Ram(read_addr, write_addr, read_clk, write_clk, we, data, q);
wire _0000_;
wire _0001_;
wire _0002_;
wire _0003_;
wire _0004_;
wire _0005_;
wire _0006_;
wire _0007_;
wire _0008_;
wire _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire _0013_;
wire _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire _0031_;
wire _0032_;
wire _0033_;
wire _0034_;
wire _0035_;
wire _0036_;
wire _0037_;
wire _0038_;
wire _0039_;
wire _0040_;
wire _0041_;
wire _0042_;
wire _0043_;
wire _0044_;
wire _0045_;
wire _0046_;
wire _0047_;
wire _0048_;
wire _0049_;
wire _0050_;
wire _0051_;
wire _0052_;
wire _0053_;
wire _0054_;
wire _0055_;
wire _0056_;
wire _0057_;
wire _0058_;
wire _0059_;
wire _0060_;
wire _0061_;
wire _0062_;
wire _0063_;
wire _0064_;
wire _0065_;
wire _0066_;
wire _0067_;
wire _0068_;
wire _0069_;
wire _0070_;
wire _0071_;
wire _0072_;
wire _0073_;
wire _0074_;
wire _0075_;
wire _0076_;
wire _0077_;
wire _0078_;
wire _0079_;
wire _0080_;
wire _0081_;
wire _0082_;
wire _0083_;
wire _0084_;
wire _0085_;
wire _0086_;
wire _0087_;
wire _0088_;
wire _0089_;
wire _0090_;
wire _0091_;
wire _0092_;
wire _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire _0144_;
wire _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire _0278_;
wire _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0327_;
wire _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire _0350_;
wire _0351_;
wire _0352_;
wire _0353_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0357_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0366_;
wire _0367_;
wire _0368_;
wire _0369_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire _0427_;
wire _0428_;
wire _0429_;
wire _0430_;
wire _0431_;
wire _0432_;
wire _0433_;
wire _0434_;
wire _0435_;
wire _0436_;
wire _0437_;
wire _0438_;
wire _0439_;
wire _0440_;
wire _0441_;
wire _0442_;
wire _0443_;
wire _0444_;
wire _0445_;
wire _0446_;
wire _0447_;
wire _0448_;
wire _0449_;
wire _0450_;
wire _0451_;
wire _0452_;
wire _0453_;
wire _0454_;
wire _0455_;
wire _0456_;
wire _0457_;
wire _0458_;
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire _0487_;
wire _0488_;
wire _0489_;
wire _0490_;
wire _0491_;
wire _0492_;
wire _0493_;
wire _0494_;
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0542_;
wire _0543_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire _0610_;
wire _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire _0616_;
wire _0617_;
wire _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire _0622_;
wire _0623_;
wire _0624_;
wire _0625_;
wire _0626_;
wire _0627_;
wire _0628_;
wire _0629_;
wire _0630_;
wire _0631_;
wire _0632_;
wire _0633_;
wire _0634_;
wire _0635_;
wire _0636_;
wire _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire _0651_;
wire _0652_;
wire _0653_;
wire _0654_;
wire _0655_;
wire _0656_;
wire _0657_;
wire _0658_;
wire _0659_;
wire _0660_;
wire _0661_;
wire _0662_;
wire _0663_;
wire _0664_;
wire _0665_;
wire _0666_;
wire _0667_;
wire _0668_;
wire _0669_;
wire _0670_;
wire _0671_;
wire _0672_;
wire _0673_;
wire _0674_;
wire _0675_;
wire _0676_;
wire _0677_;
wire _0678_;
wire _0679_;
wire _0680_;
wire _0681_;
wire _0682_;
wire _0683_;
wire _0684_;
wire _0685_;
wire _0686_;
wire _0687_;
wire _0688_;
wire _0689_;
wire _0690_;
wire _0691_;
wire _0692_;
wire _0693_;
wire _0694_;
wire _0695_;
wire _0696_;
wire _0697_;
wire _0698_;
wire _0699_;
wire _0700_;
wire _0701_;
wire _0702_;
wire _0703_;
wire _0704_;
wire _0705_;
wire _0706_;
wire _0707_;
wire _0708_;
wire _0709_;
wire _0710_;
wire _0711_;
wire _0712_;
wire _0713_;
wire _0714_;
wire _0715_;
wire _0716_;
wire _0717_;
wire _0718_;
wire _0719_;
wire _0720_;
wire _0721_;
wire _0722_;
wire _0723_;
wire _0724_;
wire _0725_;
wire _0726_;
wire _0727_;
wire _0728_;
wire _0729_;
wire _0730_;
wire _0731_;
wire _0732_;
wire _0733_;
wire _0734_;
wire _0735_;
wire _0736_;
wire _0737_;
wire _0738_;
wire _0739_;
wire _0740_;
wire _0741_;
wire _0742_;
wire _0743_;
wire _0744_;
wire _0745_;
wire _0746_;
wire _0747_;
wire _0748_;
wire _0749_;
wire _0750_;
wire _0751_;
wire _0752_;
wire _0753_;
wire _0754_;
wire _0755_;
wire _0756_;
wire _0757_;
wire _0758_;
wire _0759_;
wire _0760_;
wire _0761_;
wire _0762_;
wire _0763_;
wire _0764_;
wire _0765_;
wire _0766_;
wire _0767_;
wire _0768_;
wire _0769_;
wire _0770_;
wire _0771_;
wire _0772_;
wire _0773_;
wire _0774_;
wire _0775_;
wire _0776_;
wire _0777_;
wire _0778_;
wire _0779_;
wire _0780_;
wire _0781_;
wire _0782_;
wire _0783_;
wire _0784_;
wire _0785_;
wire _0786_;
wire _0787_;
wire _0788_;
wire _0789_;
wire _0790_;
wire _0791_;
wire _0792_;
wire _0793_;
wire _0794_;
wire _0795_;
wire _0796_;
wire _0797_;
wire _0798_;
wire _0799_;
wire _0800_;
wire _0801_;
wire _0802_;
wire _0803_;
wire _0804_;
wire _0805_;
wire _0806_;
wire _0807_;
wire _0808_;
wire _0809_;
wire _0810_;
wire _0811_;
wire _0812_;
wire _0813_;
wire _0814_;
wire _0815_;
wire _0816_;
wire _0817_;
wire _0818_;
wire _0819_;
wire _0820_;
wire _0821_;
wire _0822_;
wire _0823_;
wire _0824_;
wire _0825_;
wire _0826_;
wire _0827_;
wire _0828_;
wire _0829_;
wire _0830_;
wire _0831_;
wire _0832_;
wire _0833_;
wire _0834_;
wire _0835_;
wire _0836_;
wire _0837_;
wire _0838_;
wire _0839_;
wire _0840_;
wire _0841_;
wire _0842_;
wire _0843_;
wire _0844_;
wire _0845_;
wire _0846_;
wire _0847_;
wire _0848_;
wire _0849_;
wire _0850_;
wire _0851_;
wire _0852_;
wire _0853_;
wire _0854_;
wire _0855_;
wire _0856_;
wire _0857_;
wire _0858_;
wire _0859_;
wire _0860_;
wire _0861_;
wire _0862_;
wire _0863_;
wire _0864_;
wire _0865_;
wire _0866_;
wire _0867_;
wire _0868_;
wire _0869_;
wire _0870_;
wire _0871_;
wire _0872_;
wire _0873_;
wire _0874_;
wire _0875_;
wire _0876_;
wire _0877_;
wire _0878_;
wire _0879_;
wire _0880_;
wire _0881_;
wire _0882_;
wire _0883_;
wire _0884_;
wire _0885_;
wire _0886_;
wire _0887_;
wire _0888_;
wire _0889_;
wire _0890_;
wire _0891_;
wire _0892_;
wire _0893_;
wire _0894_;
wire _0895_;
wire _0896_;
wire _0897_;
wire _0898_;
wire _0899_;
wire _0900_;
wire _0901_;
wire _0902_;
wire _0903_;
wire _0904_;
wire _0905_;
wire _0906_;
wire _0907_;
wire _0908_;
wire _0909_;
wire _0910_;
wire _0911_;
wire _0912_;
wire _0913_;
wire _0914_;
wire _0915_;
wire _0916_;
wire _0917_;
wire _0918_;
wire _0919_;
wire _0920_;
wire _0921_;
wire _0922_;
wire _0923_;
wire _0924_;
wire _0925_;
wire _0926_;
wire _0927_;
wire _0928_;
wire _0929_;
wire _0930_;
wire _0931_;
wire _0932_;
wire _0933_;
wire _0934_;
wire _0935_;
wire _0936_;
wire _0937_;
wire _0938_;
wire _0939_;
wire _0940_;
wire _0941_;
wire _0942_;
wire _0943_;
wire _0944_;
wire _0945_;
wire _0946_;
wire _0947_;
wire _0948_;
wire _0949_;
wire _0950_;
wire _0951_;
wire _0952_;
wire _0953_;
wire _0954_;
wire _0955_;
wire _0956_;
wire _0957_;
wire _0958_;
wire _0959_;
wire _0960_;
wire _0961_;
wire _0962_;
wire _0963_;
wire _0964_;
wire _0965_;
wire _0966_;
wire _0967_;
wire _0968_;
wire _0969_;
wire _0970_;
wire _0971_;
wire _0972_;
wire _0973_;
wire _0974_;
wire _0975_;
wire _0976_;
wire _0977_;
wire _0978_;
wire _0979_;
wire _0980_;
wire _0981_;
wire _0982_;
wire _0983_;
wire _0984_;
wire _0985_;
wire _0986_;
wire _0987_;
wire _0988_;
wire _0989_;
wire _0990_;
wire _0991_;
wire _0992_;
wire _0993_;
wire _0994_;
wire _0995_;
wire _0996_;
wire _0997_;
wire _0998_;
wire _0999_;
wire _1000_;
wire _1001_;
wire _1002_;
wire _1003_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1023_;
wire _1024_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1033_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1130_;
wire _1131_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1138_;
wire _1139_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1151_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1161_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire _1218_;
wire _1219_;
wire _1220_;
wire _1221_;
wire _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire _1227_;
wire _1228_;
wire _1229_;
wire _1230_;
wire _1231_;
wire _1232_;
wire _1233_;
wire _1234_;
wire _1235_;
wire _1236_;
wire _1237_;
wire _1238_;
wire _1239_;
wire _1240_;
wire _1241_;
wire _1242_;
wire _1243_;
wire _1244_;
wire _1245_;
wire _1246_;
wire _1247_;
wire _1248_;
wire _1249_;
wire _1250_;
wire _1251_;
wire _1252_;
wire _1253_;
wire _1254_;
wire _1255_;
wire _1256_;
wire _1257_;
wire _1258_;
wire _1259_;
wire _1260_;
wire _1261_;
wire _1262_;
wire _1263_;
wire _1264_;
wire _1265_;
wire _1266_;
wire _1267_;
wire _1268_;
wire _1269_;
wire _1270_;
wire _1271_;
wire _1272_;
wire _1273_;
wire _1274_;
wire _1275_;
wire _1276_;
wire _1277_;
wire _1278_;
wire _1279_;
wire _1280_;
wire _1281_;
wire _1282_;
wire _1283_;
wire _1284_;
wire _1285_;
wire _1286_;
wire _1287_;
wire _1288_;
wire _1289_;
wire _1290_;
wire _1291_;
wire _1292_;
wire _1293_;
wire _1294_;
wire _1295_;
wire _1296_;
wire _1297_;
wire _1298_;
wire _1299_;
wire _1300_;
wire _1301_;
wire _1302_;
wire _1303_;
wire _1304_;
wire _1305_;
wire _1306_;
wire _1307_;
wire _1308_;
wire _1309_;
wire _1310_;
wire _1311_;
wire _1312_;
wire _1313_;
wire _1314_;
wire _1315_;
wire _1316_;
wire _1317_;
wire _1318_;
wire _1319_;
wire _1320_;
wire _1321_;
wire _1322_;
wire _1323_;
wire _1324_;
wire _1325_;
wire _1326_;
wire _1327_;
wire _1328_;
wire _1329_;
wire _1330_;
wire _1331_;
wire _1332_;
wire _1333_;
wire _1334_;
wire _1335_;
wire _1336_;
wire _1337_;
wire _1338_;
wire _1339_;
wire _1340_;
wire _1341_;
wire _1342_;
wire _1343_;
wire _1344_;
wire _1345_;
wire _1346_;
wire _1347_;
wire _1348_;
wire _1349_;
wire _1350_;
wire _1351_;
wire _1352_;
wire _1353_;
wire _1354_;
wire _1355_;
wire _1356_;
wire _1357_;
wire _1358_;
wire _1359_;
wire _1360_;
wire _1361_;
wire _1362_;
wire _1363_;
wire _1364_;
wire _1365_;
wire _1366_;
wire _1367_;
wire _1368_;
wire _1369_;
wire _1370_;
wire _1371_;
wire _1372_;
wire _1373_;
wire _1374_;
wire _1375_;
wire _1376_;
wire _1377_;
wire _1378_;
wire _1379_;
wire _1380_;
wire _1381_;
wire _1382_;
wire _1383_;
wire _1384_;
wire _1385_;
wire _1386_;
wire _1387_;
wire _1388_;
wire _1389_;
wire _1390_;
wire _1391_;
wire _1392_;
wire _1393_;
wire _1394_;
wire _1395_;
wire _1396_;
wire _1397_;
wire _1398_;
wire _1399_;
wire _1400_;
wire _1401_;
wire _1402_;
wire _1403_;
wire _1404_;
wire _1405_;
wire _1406_;
wire _1407_;
wire _1408_;
wire _1409_;
wire _1410_;
wire _1411_;
wire _1412_;
wire _1413_;
wire _1414_;
wire _1415_;
wire _1416_;
wire _1417_;
wire _1418_;
wire _1419_;
wire _1420_;
wire _1421_;
wire _1422_;
wire _1423_;
wire _1424_;
wire _1425_;
wire _1426_;
wire _1427_;
wire _1428_;
wire _1429_;
wire _1430_;
wire _1431_;
wire _1432_;
wire _1433_;
wire _1434_;
wire _1435_;
wire _1436_;
wire _1437_;
wire _1438_;
wire _1439_;
wire _1440_;
wire _1441_;
wire _1442_;
wire _1443_;
wire _1444_;
wire _1445_;
wire _1446_;
wire _1447_;
wire _1448_;
wire _1449_;
wire _1450_;
wire _1451_;
wire _1452_;
wire _1453_;
wire _1454_;
wire _1455_;
wire _1456_;
wire _1457_;
wire _1458_;
wire _1459_;
wire _1460_;
wire _1461_;
wire _1462_;
wire _1463_;
wire _1464_;
wire _1465_;
wire _1466_;
wire _1467_;
wire _1468_;
wire _1469_;
wire _1470_;
wire _1471_;
wire _1472_;
wire _1473_;
wire _1474_;
wire _1475_;
wire _1476_;
wire _1477_;
wire _1478_;
wire _1479_;
wire _1480_;
wire _1481_;
wire _1482_;
wire _1483_;
wire _1484_;
wire _1485_;
wire _1486_;
wire _1487_;
wire _1488_;
wire _1489_;
wire _1490_;
wire _1491_;
wire _1492_;
wire _1493_;
wire _1494_;
wire _1495_;
wire _1496_;
wire _1497_;
wire _1498_;
wire _1499_;
wire _1500_;
wire _1501_;
wire _1502_;
wire _1503_;
wire _1504_;
wire _1505_;
wire _1506_;
wire _1507_;
wire _1508_;
wire _1509_;
wire _1510_;
wire _1511_;
wire _1512_;
wire _1513_;
wire _1514_;
wire _1515_;
wire _1516_;
wire _1517_;
wire _1518_;
wire _1519_;
wire _1520_;
wire _1521_;
wire _1522_;
wire _1523_;
wire _1524_;
wire _1525_;
wire _1526_;
wire _1527_;
wire _1528_;
wire _1529_;
wire _1530_;
wire _1531_;
wire _1532_;
wire _1533_;
wire _1534_;
wire _1535_;
wire _1536_;
wire _1537_;
wire _1538_;
wire _1539_;
wire _1540_;
wire _1541_;
wire _1542_;
wire _1543_;
wire _1544_;
wire _1545_;
wire _1546_;
wire _1547_;
wire _1548_;
wire _1549_;
wire _1550_;
wire _1551_;
wire _1552_;
wire _1553_;
wire _1554_;
wire _1555_;
wire _1556_;
wire _1557_;
wire _1558_;
wire _1559_;
wire _1560_;
wire _1561_;
wire _1562_;
wire _1563_;
wire _1564_;
wire _1565_;
wire _1566_;
wire _1567_;
wire _1568_;
wire _1569_;
wire _1570_;
wire _1571_;
wire _1572_;
wire _1573_;
wire _1574_;
wire _1575_;
wire _1576_;
wire _1577_;
wire _1578_;
wire _1579_;
wire _1580_;
wire _1581_;
wire _1582_;
wire _1583_;
wire _1584_;
wire _1585_;
wire _1586_;
wire _1587_;
wire _1588_;
wire _1589_;
wire _1590_;
wire _1591_;
wire _1592_;
wire _1593_;
wire _1594_;
wire _1595_;
wire _1596_;
wire _1597_;
wire _1598_;
wire _1599_;
wire _1600_;
wire _1601_;
wire _1602_;
wire _1603_;
wire _1604_;
wire _1605_;
wire _1606_;
wire _1607_;
wire _1608_;
wire _1609_;
wire _1610_;
wire _1611_;
wire _1612_;
wire _1613_;
wire _1614_;
wire _1615_;
wire _1616_;
wire _1617_;
wire _1618_;
wire _1619_;
wire _1620_;
wire _1621_;
wire _1622_;
wire _1623_;
wire _1624_;
wire _1625_;
wire _1626_;
wire _1627_;
wire _1628_;
wire _1629_;
wire _1630_;
input [15:0] data;
wire [15:0] \mem[0] ;
wire [15:0] \mem[10] ;
wire [15:0] \mem[11] ;
wire [15:0] \mem[12] ;
wire [15:0] \mem[13] ;
wire [15:0] \mem[14] ;
wire [15:0] \mem[15] ;
wire [15:0] \mem[1] ;
wire [15:0] \mem[2] ;
wire [15:0] \mem[3] ;
wire [15:0] \mem[4] ;
wire [15:0] \mem[5] ;
wire [15:0] \mem[6] ;
wire [15:0] \mem[7] ;
wire [15:0] \mem[8] ;
wire [15:0] \mem[9] ;
output [15:0] q;
input [3:0] read_addr;
input read_clk;
input we;
input [3:0] write_addr;
input write_clk;
NOT _1631_ (.A(\mem[14] [0]),.Y(_1279_));
NOT _1632_ (.A(\mem[14] [1]),.Y(_1280_));
NOT _1633_ (.A(\mem[14] [3]),.Y(_1281_));
NOT _1634_ (.A(\mem[14] [4]),.Y(_1282_));
NOT _1635_ (.A(\mem[14] [5]),.Y(_1283_));
NOT _1636_ (.A(\mem[14] [6]),.Y(_1284_));
NOT _1637_ (.A(\mem[14] [7]),.Y(_1285_));
NOT _1638_ (.A(\mem[14] [8]),.Y(_1286_));
NOT _1639_ (.A(\mem[14] [9]),.Y(_1287_));
NOT _1640_ (.A(\mem[14] [10]),.Y(_1288_));
NOT _1641_ (.A(\mem[14] [11]),.Y(_1289_));
NOT _1642_ (.A(\mem[14] [12]),.Y(_1290_));
NOT _1643_ (.A(\mem[14] [13]),.Y(_1291_));
NOT _1644_ (.A(\mem[14] [14]),.Y(_1292_));
NOT _1645_ (.A(\mem[14] [15]),.Y(_1293_));
NOT _1646_ (.A(\mem[15] [0]),.Y(_1294_));
NOT _1647_ (.A(\mem[15] [1]),.Y(_1295_));
NOT _1648_ (.A(\mem[15] [3]),.Y(_1296_));
NOT _1649_ (.A(\mem[15] [4]),.Y(_1297_));
NOT _1650_ (.A(\mem[15] [5]),.Y(_1298_));
NOT _1651_ (.A(\mem[15] [6]),.Y(_1299_));
NOT _1652_ (.A(\mem[15] [7]),.Y(_1300_));
NOT _1653_ (.A(\mem[15] [8]),.Y(_1301_));
NOT _1654_ (.A(\mem[15] [9]),.Y(_1302_));
NOT _1655_ (.A(\mem[15] [10]),.Y(_1303_));
NOT _1656_ (.A(\mem[15] [11]),.Y(_1304_));
NOT _1657_ (.A(\mem[15] [12]),.Y(_1305_));
NOT _1658_ (.A(\mem[15] [13]),.Y(_1306_));
NOT _1659_ (.A(\mem[15] [14]),.Y(_1307_));
NOT _1660_ (.A(\mem[15] [15]),.Y(_1308_));
NOT _1661_ (.A(write_addr[0]),.Y(_1309_));
NOT _1662_ (.A(we),.Y(_1310_));
NOT _1663_ (.A(write_addr[1]),.Y(_1311_));
NOT _1664_ (.A(write_addr[2]),.Y(_1312_));
NOT _1665_ (.A(write_addr[3]),.Y(_1313_));
NOT _1666_ (.A(data[0]),.Y(_1314_));
NOT _1667_ (.A(data[1]),.Y(_1315_));
NOT _1668_ (.A(data[2]),.Y(_1316_));
NOT _1669_ (.A(data[3]),.Y(_1317_));
NOT _1670_ (.A(data[4]),.Y(_1318_));
NOT _1671_ (.A(data[5]),.Y(_1319_));
NOT _1672_ (.A(data[6]),.Y(_1320_));
NOT _1673_ (.A(data[7]),.Y(_1321_));
NOT _1674_ (.A(data[8]),.Y(_1322_));
NOT _1675_ (.A(data[9]),.Y(_1323_));
NOT _1676_ (.A(data[10]),.Y(_1324_));
NOT _1677_ (.A(data[11]),.Y(_1325_));
NOT _1678_ (.A(data[12]),.Y(_1326_));
NOT _1679_ (.A(data[13]),.Y(_1327_));
NOT _1680_ (.A(data[14]),.Y(_1328_));
NOT _1681_ (.A(data[15]),.Y(_1329_));
NOT _1682_ (.A(read_addr[3]),.Y(_1330_));
NOT _1683_ (.A(read_addr[2]),.Y(_1331_));
NOT _1684_ (.A(read_addr[1]),.Y(_1332_));
NOT _1685_ (.A(read_addr[0]),.Y(_1333_));
NOT _1686_ (.A(\mem[3] [0]),.Y(_1334_));
NOT _1687_ (.A(\mem[3] [1]),.Y(_1335_));
NOT _1688_ (.A(\mem[3] [9]),.Y(_1336_));
NOT _1689_ (.A(\mem[3] [10]),.Y(_1337_));
NOT _1690_ (.A(\mem[3] [14]),.Y(_1338_));
NOT _1691_ (.A(\mem[8] [3]),.Y(_1339_));
NOT _1692_ (.A(\mem[9] [3]),.Y(_1340_));
NOT _1693_ (.A(\mem[8] [5]),.Y(_1341_));
NOT _1694_ (.A(\mem[9] [5]),.Y(_1342_));
NOT _1695_ (.A(\mem[8] [7]),.Y(_1343_));
NOT _1696_ (.A(\mem[9] [7]),.Y(_1344_));
NOT _1697_ (.A(\mem[8] [15]),.Y(_1345_));
NOT _1698_ (.A(\mem[9] [15]),.Y(_1346_));
NOR _1699_ (.A(_1310_),.B(_1311_),.Y(_1347_));
NAND _1700_ (.A(we),.B(write_addr[1]),.Y(_1348_));
NOR _1701_ (.A(write_addr[0]),.B(_1348_),.Y(_1349_));
NAND _1702_ (.A(_1309_),.B(_1347_),.Y(_1350_));
NOR _1703_ (.A(_1310_),.B(_1313_),.Y(_1351_));
NAND _1704_ (.A(we),.B(write_addr[3]),.Y(_1352_));
NOR _1705_ (.A(write_addr[2]),.B(_1352_),.Y(_1353_));
NAND _1706_ (.A(_1312_),.B(_1351_),.Y(_1354_));
NOR _1707_ (.A(_1350_),.B(_1354_),.Y(_1355_));
NAND _1708_ (.A(_1349_),.B(_1353_),.Y(_1356_));
NOR _1709_ (.A(_1310_),.B(_1317_),.Y(_1357_));
NAND _1710_ (.A(_1355_),.B(_1357_),.Y(_1358_));
NAND _1711_ (.A(\mem[10] [3]),.B(_1356_),.Y(_1359_));
NAND _1712_ (.A(_1358_),.B(_1359_),.Y(_0041_));
NAND _1713_ (.A(\mem[10] [4]),.B(_1356_),.Y(_1360_));
NOR _1714_ (.A(_1310_),.B(_1318_),.Y(_1361_));
NAND _1715_ (.A(_1355_),.B(_1361_),.Y(_1362_));
NAND _1716_ (.A(_1360_),.B(_1362_),.Y(_0042_));
NAND _1717_ (.A(\mem[10] [5]),.B(_1356_),.Y(_1363_));
NOR _1718_ (.A(_1310_),.B(_1319_),.Y(_1364_));
NAND _1719_ (.A(_1355_),.B(_1364_),.Y(_1365_));
NAND _1720_ (.A(_1363_),.B(_1365_),.Y(_0043_));
NAND _1721_ (.A(\mem[10] [6]),.B(_1356_),.Y(_1366_));
NOR _1722_ (.A(_1310_),.B(_1320_),.Y(_1367_));
NAND _1723_ (.A(_1355_),.B(_1367_),.Y(_1368_));
NAND _1724_ (.A(_1366_),.B(_1368_),.Y(_0044_));
NAND _1725_ (.A(\mem[10] [7]),.B(_1356_),.Y(_1369_));
NOR _1726_ (.A(_1310_),.B(_1321_),.Y(_1370_));
NAND _1727_ (.A(_1355_),.B(_1370_),.Y(_1371_));
NAND _1728_ (.A(_1369_),.B(_1371_),.Y(_0045_));
NOR _1729_ (.A(_1310_),.B(_1322_),.Y(_1372_));
NAND _1730_ (.A(_1355_),.B(_1372_),.Y(_1373_));
NAND _1731_ (.A(\mem[10] [8]),.B(_1356_),.Y(_1374_));
NAND _1732_ (.A(_1373_),.B(_1374_),.Y(_0046_));
NOR _1733_ (.A(_1310_),.B(_1323_),.Y(_1375_));
NAND _1734_ (.A(_1355_),.B(_1375_),.Y(_1376_));
NAND _1735_ (.A(\mem[10] [9]),.B(_1356_),.Y(_1377_));
NAND _1736_ (.A(_1376_),.B(_1377_),.Y(_0047_));
NAND _1737_ (.A(\mem[10] [10]),.B(_1356_),.Y(_1378_));
NOR _1738_ (.A(_1310_),.B(_1324_),.Y(_1379_));
NAND _1739_ (.A(_1355_),.B(_1379_),.Y(_1380_));
NAND _1740_ (.A(_1378_),.B(_1380_),.Y(_0033_));
NAND _1741_ (.A(\mem[10] [11]),.B(_1356_),.Y(_1381_));
NOR _1742_ (.A(_1310_),.B(_1325_),.Y(_1382_));
NAND _1743_ (.A(_1355_),.B(_1382_),.Y(_1383_));
NAND _1744_ (.A(_1381_),.B(_1383_),.Y(_0034_));
NAND _1745_ (.A(\mem[10] [12]),.B(_1356_),.Y(_1384_));
NOR _1746_ (.A(_1310_),.B(_1326_),.Y(_1385_));
NAND _1747_ (.A(_1355_),.B(_1385_),.Y(_1386_));
NAND _1748_ (.A(_1384_),.B(_1386_),.Y(_0035_));
NAND _1749_ (.A(\mem[10] [13]),.B(_1356_),.Y(_1387_));
NOR _1750_ (.A(_1310_),.B(_1327_),.Y(_1388_));
NAND _1751_ (.A(_1355_),.B(_1388_),.Y(_1389_));
NAND _1752_ (.A(_1387_),.B(_1389_),.Y(_0036_));
NAND _1753_ (.A(\mem[10] [14]),.B(_1356_),.Y(_1390_));
NOR _1754_ (.A(_1310_),.B(_1328_),.Y(_1391_));
NAND _1755_ (.A(_1355_),.B(_1391_),.Y(_1392_));
NAND _1756_ (.A(_1390_),.B(_1392_),.Y(_0037_));
NOR _1757_ (.A(_1310_),.B(_1329_),.Y(_1393_));
NAND _1758_ (.A(_1355_),.B(_1393_),.Y(_1394_));
NAND _1759_ (.A(\mem[10] [15]),.B(_1356_),.Y(_1395_));
NAND _1760_ (.A(_1394_),.B(_1395_),.Y(_0038_));
NOR _1761_ (.A(_1309_),.B(_1310_),.Y(_1396_));
NAND _1762_ (.A(write_addr[0]),.B(we),.Y(_1397_));
NOR _1763_ (.A(_1309_),.B(_1348_),.Y(_1398_));
NAND _1764_ (.A(write_addr[0]),.B(_1347_),.Y(_1399_));
NOR _1765_ (.A(_1354_),.B(_1399_),.Y(_1400_));
NAND _1766_ (.A(_1353_),.B(_1398_),.Y(_1401_));
NOR _1767_ (.A(_1310_),.B(_1314_),.Y(_1402_));
NAND _1768_ (.A(_1400_),.B(_1402_),.Y(_1403_));
NAND _1769_ (.A(\mem[11] [0]),.B(_1401_),.Y(_1404_));
NAND _1770_ (.A(_1403_),.B(_1404_),.Y(_0048_));
NOR _1771_ (.A(_1310_),.B(_1315_),.Y(_1405_));
NAND _1772_ (.A(_1400_),.B(_1405_),.Y(_1406_));
NAND _1773_ (.A(\mem[11] [1]),.B(_1401_),.Y(_1407_));
NAND _1774_ (.A(_1406_),.B(_1407_),.Y(_0055_));
NOR _1775_ (.A(_1310_),.B(_1316_),.Y(_1408_));
NAND _1776_ (.A(_1400_),.B(_1408_),.Y(_1409_));
NAND _1777_ (.A(\mem[11] [2]),.B(_1401_),.Y(_1410_));
NAND _1778_ (.A(_1409_),.B(_1410_),.Y(_0056_));
NAND _1779_ (.A(_1357_),.B(_1400_),.Y(_1411_));
NAND _1780_ (.A(\mem[11] [3]),.B(_1401_),.Y(_1412_));
NAND _1781_ (.A(_1411_),.B(_1412_),.Y(_0057_));
NAND _1782_ (.A(_1361_),.B(_1400_),.Y(_1413_));
NAND _1783_ (.A(\mem[11] [4]),.B(_1401_),.Y(_1414_));
NAND _1784_ (.A(_1413_),.B(_1414_),.Y(_0058_));
NAND _1785_ (.A(_1364_),.B(_1400_),.Y(_1415_));
NAND _1786_ (.A(\mem[11] [5]),.B(_1401_),.Y(_1416_));
NAND _1787_ (.A(_1415_),.B(_1416_),.Y(_0059_));
NAND _1788_ (.A(_1367_),.B(_1400_),.Y(_1417_));
NAND _1789_ (.A(\mem[11] [6]),.B(_1401_),.Y(_1418_));
NAND _1790_ (.A(_1417_),.B(_1418_),.Y(_0060_));
NAND _1791_ (.A(_1370_),.B(_1400_),.Y(_1419_));
NAND _1792_ (.A(\mem[11] [7]),.B(_1401_),.Y(_1420_));
NAND _1793_ (.A(_1419_),.B(_1420_),.Y(_0061_));
NAND _1794_ (.A(_1372_),.B(_1400_),.Y(_1421_));
NAND _1795_ (.A(\mem[11] [8]),.B(_1401_),.Y(_1422_));
NAND _1796_ (.A(_1421_),.B(_1422_),.Y(_0062_));
NAND _1797_ (.A(_1375_),.B(_1400_),.Y(_1423_));
NAND _1798_ (.A(\mem[11] [9]),.B(_1401_),.Y(_1424_));
NAND _1799_ (.A(_1423_),.B(_1424_),.Y(_0063_));
NAND _1800_ (.A(_1379_),.B(_1400_),.Y(_1425_));
NAND _1801_ (.A(\mem[11] [10]),.B(_1401_),.Y(_1426_));
NAND _1802_ (.A(_1425_),.B(_1426_),.Y(_0049_));
NAND _1803_ (.A(_1382_),.B(_1400_),.Y(_1427_));
NAND _1804_ (.A(\mem[11] [11]),.B(_1401_),.Y(_1428_));
NAND _1805_ (.A(_1427_),.B(_1428_),.Y(_0050_));
NAND _1806_ (.A(_1385_),.B(_1400_),.Y(_1429_));
NAND _1807_ (.A(\mem[11] [12]),.B(_1401_),.Y(_1430_));
NAND _1808_ (.A(_1429_),.B(_1430_),.Y(_0051_));
NAND _1809_ (.A(_1388_),.B(_1400_),.Y(_1431_));
NAND _1810_ (.A(\mem[11] [13]),.B(_1401_),.Y(_1432_));
NAND _1811_ (.A(_1431_),.B(_1432_),.Y(_0052_));
NAND _1812_ (.A(_1391_),.B(_1400_),.Y(_1433_));
NAND _1813_ (.A(\mem[11] [14]),.B(_1401_),.Y(_1434_));
NAND _1814_ (.A(_1433_),.B(_1434_),.Y(_0053_));
NAND _1815_ (.A(_1393_),.B(_1400_),.Y(_1435_));
NAND _1816_ (.A(\mem[11] [15]),.B(_1401_),.Y(_1436_));
NAND _1817_ (.A(_1435_),.B(_1436_),.Y(_0054_));
NOR _1818_ (.A(_1347_),.B(_1396_),.Y(_1437_));
NAND _1819_ (.A(_1348_),.B(_1397_),.Y(_1438_));
NOR _1820_ (.A(_1310_),.B(_1312_),.Y(_1439_));
NAND _1821_ (.A(we),.B(write_addr[2]),.Y(_1440_));
NOR _1822_ (.A(_1313_),.B(_1440_),.Y(_1441_));
NAND _1823_ (.A(write_addr[3]),.B(_1439_),.Y(_1442_));
NOR _1824_ (.A(_1438_),.B(_1442_),.Y(_1443_));
NAND _1825_ (.A(_1437_),.B(_1441_),.Y(_1444_));
NAND _1826_ (.A(_1402_),.B(_1443_),.Y(_1445_));
NAND _1827_ (.A(\mem[12] [0]),.B(_1444_),.Y(_1446_));
NAND _1828_ (.A(_1445_),.B(_1446_),.Y(_0064_));
NAND _1829_ (.A(_1405_),.B(_1443_),.Y(_1447_));
NAND _1830_ (.A(\mem[12] [1]),.B(_1444_),.Y(_1448_));
NAND _1831_ (.A(_1447_),.B(_1448_),.Y(_0071_));
NAND _1832_ (.A(_1408_),.B(_1443_),.Y(_1449_));
NAND _1833_ (.A(\mem[12] [2]),.B(_1444_),.Y(_1450_));
NAND _1834_ (.A(_1449_),.B(_1450_),.Y(_0072_));
NAND _1835_ (.A(_1357_),.B(_1443_),.Y(_1451_));
NAND _1836_ (.A(\mem[12] [3]),.B(_1444_),.Y(_1452_));
NAND _1837_ (.A(_1451_),.B(_1452_),.Y(_0073_));
NAND _1838_ (.A(_1361_),.B(_1443_),.Y(_1453_));
NAND _1839_ (.A(\mem[12] [4]),.B(_1444_),.Y(_1454_));
NAND _1840_ (.A(_1453_),.B(_1454_),.Y(_0074_));
NAND _1841_ (.A(_1364_),.B(_1443_),.Y(_1455_));
NAND _1842_ (.A(\mem[12] [5]),.B(_1444_),.Y(_1456_));
NAND _1843_ (.A(_1455_),.B(_1456_),.Y(_0075_));
NAND _1844_ (.A(_1367_),.B(_1443_),.Y(_1457_));
NAND _1845_ (.A(\mem[12] [6]),.B(_1444_),.Y(_1458_));
NAND _1846_ (.A(_1457_),.B(_1458_),.Y(_0076_));
NAND _1847_ (.A(_1370_),.B(_1443_),.Y(_1459_));
NAND _1848_ (.A(\mem[12] [7]),.B(_1444_),.Y(_1460_));
NAND _1849_ (.A(_1459_),.B(_1460_),.Y(_0077_));
NAND _1850_ (.A(_1372_),.B(_1443_),.Y(_1461_));
NAND _1851_ (.A(\mem[12] [8]),.B(_1444_),.Y(_1462_));
NAND _1852_ (.A(_1461_),.B(_1462_),.Y(_0078_));
NAND _1853_ (.A(_1375_),.B(_1443_),.Y(_1463_));
NAND _1854_ (.A(\mem[12] [9]),.B(_1444_),.Y(_1464_));
NAND _1855_ (.A(_1463_),.B(_1464_),.Y(_0079_));
NAND _1856_ (.A(_1379_),.B(_1443_),.Y(_1465_));
NAND _1857_ (.A(\mem[12] [10]),.B(_1444_),.Y(_1466_));
NAND _1858_ (.A(_1465_),.B(_1466_),.Y(_0065_));
NAND _1859_ (.A(_1382_),.B(_1443_),.Y(_1467_));
NAND _1860_ (.A(\mem[12] [11]),.B(_1444_),.Y(_1468_));
NAND _1861_ (.A(_1467_),.B(_1468_),.Y(_0066_));
NAND _1862_ (.A(_1385_),.B(_1443_),.Y(_1469_));
NAND _1863_ (.A(\mem[12] [12]),.B(_1444_),.Y(_1470_));
NAND _1864_ (.A(_1469_),.B(_1470_),.Y(_0067_));
NAND _1865_ (.A(_1388_),.B(_1443_),.Y(_1471_));
NAND _1866_ (.A(\mem[12] [13]),.B(_1444_),.Y(_1472_));
NAND _1867_ (.A(_1471_),.B(_1472_),.Y(_0068_));
NAND _1868_ (.A(_1391_),.B(_1443_),.Y(_1473_));
NAND _1869_ (.A(\mem[12] [14]),.B(_1444_),.Y(_1474_));
NAND _1870_ (.A(_1473_),.B(_1474_),.Y(_0069_));
NAND _1871_ (.A(_1393_),.B(_1443_),.Y(_1475_));
NAND _1872_ (.A(\mem[12] [15]),.B(_1444_),.Y(_1476_));
NAND _1873_ (.A(_1475_),.B(_1476_),.Y(_0070_));
NOR _1874_ (.A(write_addr[1]),.B(_1397_),.Y(_1477_));
NAND _1875_ (.A(_1311_),.B(_1396_),.Y(_1478_));
NOR _1876_ (.A(_1442_),.B(_1478_),.Y(_1479_));
NAND _1877_ (.A(_1441_),.B(_1477_),.Y(_1480_));
NAND _1878_ (.A(_1402_),.B(_1479_),.Y(_1481_));
NAND _1879_ (.A(\mem[13] [0]),.B(_1480_),.Y(_1482_));
NAND _1880_ (.A(_1481_),.B(_1482_),.Y(_0080_));
NAND _1881_ (.A(_1405_),.B(_1479_),.Y(_1483_));
NAND _1882_ (.A(\mem[13] [1]),.B(_1480_),.Y(_1484_));
NAND _1883_ (.A(_1483_),.B(_1484_),.Y(_0087_));
NAND _1884_ (.A(_1408_),.B(_1479_),.Y(_1485_));
NAND _1885_ (.A(\mem[13] [2]),.B(_1480_),.Y(_1486_));
NAND _1886_ (.A(_1485_),.B(_1486_),.Y(_0088_));
NAND _1887_ (.A(_1357_),.B(_1479_),.Y(_1487_));
NAND _1888_ (.A(\mem[13] [3]),.B(_1480_),.Y(_1488_));
NAND _1889_ (.A(_1487_),.B(_1488_),.Y(_0089_));
NAND _1890_ (.A(_1361_),.B(_1479_),.Y(_1489_));
NAND _1891_ (.A(\mem[13] [4]),.B(_1480_),.Y(_1490_));
NAND _1892_ (.A(_1489_),.B(_1490_),.Y(_0090_));
NAND _1893_ (.A(_1364_),.B(_1479_),.Y(_1491_));
NAND _1894_ (.A(\mem[13] [5]),.B(_1480_),.Y(_1492_));
NAND _1895_ (.A(_1491_),.B(_1492_),.Y(_0091_));
NAND _1896_ (.A(_1367_),.B(_1479_),.Y(_1493_));
NAND _1897_ (.A(\mem[13] [6]),.B(_1480_),.Y(_1494_));
NAND _1898_ (.A(_1493_),.B(_1494_),.Y(_0092_));
NAND _1899_ (.A(_1370_),.B(_1479_),.Y(_1495_));
NAND _1900_ (.A(\mem[13] [7]),.B(_1480_),.Y(_1496_));
NAND _1901_ (.A(_1495_),.B(_1496_),.Y(_0093_));
NAND _1902_ (.A(_1372_),.B(_1479_),.Y(_1497_));
NAND _1903_ (.A(\mem[13] [8]),.B(_1480_),.Y(_1498_));
NAND _1904_ (.A(_1497_),.B(_1498_),.Y(_0094_));
NAND _1905_ (.A(_1375_),.B(_1479_),.Y(_1499_));
NAND _1906_ (.A(\mem[13] [9]),.B(_1480_),.Y(_1500_));
NAND _1907_ (.A(_1499_),.B(_1500_),.Y(_0095_));
NAND _1908_ (.A(_1379_),.B(_1479_),.Y(_1501_));
NAND _1909_ (.A(\mem[13] [10]),.B(_1480_),.Y(_1502_));
NAND _1910_ (.A(_1501_),.B(_1502_),.Y(_0081_));
NAND _1911_ (.A(_1382_),.B(_1479_),.Y(_1503_));
NAND _1912_ (.A(\mem[13] [11]),.B(_1480_),.Y(_1504_));
NAND _1913_ (.A(_1503_),.B(_1504_),.Y(_0082_));
NAND _1914_ (.A(_1385_),.B(_1479_),.Y(_1505_));
NAND _1915_ (.A(\mem[13] [12]),.B(_1480_),.Y(_1506_));
NAND _1916_ (.A(_1505_),.B(_1506_),.Y(_0083_));
NAND _1917_ (.A(_1388_),.B(_1479_),.Y(_1507_));
NAND _1918_ (.A(\mem[13] [13]),.B(_1480_),.Y(_1508_));
NAND _1919_ (.A(_1507_),.B(_1508_),.Y(_0084_));
NAND _1920_ (.A(_1391_),.B(_1479_),.Y(_1509_));
NAND _1921_ (.A(\mem[13] [14]),.B(_1480_),.Y(_1510_));
NAND _1922_ (.A(_1509_),.B(_1510_),.Y(_0085_));
NAND _1923_ (.A(_1393_),.B(_1479_),.Y(_1511_));
NAND _1924_ (.A(\mem[13] [15]),.B(_1480_),.Y(_1512_));
NAND _1925_ (.A(_1511_),.B(_1512_),.Y(_0086_));
NOR _1926_ (.A(_1350_),.B(_1442_),.Y(_1513_));
NAND _1927_ (.A(_1349_),.B(_1441_),.Y(_1514_));
NAND _1928_ (.A(_1402_),.B(_1513_),.Y(_1515_));
NAND _1929_ (.A(\mem[14] [0]),.B(_1514_),.Y(_1516_));
NAND _1930_ (.A(_1515_),.B(_1516_),.Y(_0096_));
NAND _1931_ (.A(_1405_),.B(_1513_),.Y(_1517_));
NAND _1932_ (.A(\mem[14] [1]),.B(_1514_),.Y(_1518_));
NAND _1933_ (.A(_1517_),.B(_1518_),.Y(_0103_));
NAND _1934_ (.A(_1408_),.B(_1513_),.Y(_1519_));
NAND _1935_ (.A(\mem[14] [2]),.B(_1514_),.Y(_1520_));
NAND _1936_ (.A(_1519_),.B(_1520_),.Y(_0104_));
NAND _1937_ (.A(_1357_),.B(_1513_),.Y(_1521_));
NAND _1938_ (.A(\mem[14] [3]),.B(_1514_),.Y(_1522_));
NAND _1939_ (.A(_1521_),.B(_1522_),.Y(_0105_));
NAND _1940_ (.A(_1361_),.B(_1513_),.Y(_1523_));
NAND _1941_ (.A(\mem[14] [4]),.B(_1514_),.Y(_1524_));
NAND _1942_ (.A(_1523_),.B(_1524_),.Y(_0106_));
NAND _1943_ (.A(_1364_),.B(_1513_),.Y(_1525_));
NAND _1944_ (.A(\mem[14] [5]),.B(_1514_),.Y(_1526_));
NAND _1945_ (.A(_1525_),.B(_1526_),.Y(_0107_));
NAND _1946_ (.A(_1367_),.B(_1513_),.Y(_1527_));
NAND _1947_ (.A(\mem[14] [6]),.B(_1514_),.Y(_1528_));
NAND _1948_ (.A(_1527_),.B(_1528_),.Y(_0108_));
NAND _1949_ (.A(_1370_),.B(_1513_),.Y(_1529_));
NAND _1950_ (.A(\mem[14] [7]),.B(_1514_),.Y(_1530_));
NAND _1951_ (.A(_1529_),.B(_1530_),.Y(_0109_));
NAND _1952_ (.A(_1372_),.B(_1513_),.Y(_1531_));
NAND _1953_ (.A(\mem[14] [8]),.B(_1514_),.Y(_1532_));
NAND _1954_ (.A(_1531_),.B(_1532_),.Y(_0110_));
NAND _1955_ (.A(_1375_),.B(_1513_),.Y(_1533_));
NAND _1956_ (.A(\mem[14] [9]),.B(_1514_),.Y(_1534_));
NAND _1957_ (.A(_1533_),.B(_1534_),.Y(_0111_));
NAND _1958_ (.A(_1379_),.B(_1513_),.Y(_1535_));
NAND _1959_ (.A(\mem[14] [10]),.B(_1514_),.Y(_1536_));
NAND _1960_ (.A(_1535_),.B(_1536_),.Y(_0097_));
NAND _1961_ (.A(_1382_),.B(_1513_),.Y(_1537_));
NAND _1962_ (.A(\mem[14] [11]),.B(_1514_),.Y(_1538_));
NAND _1963_ (.A(_1537_),.B(_1538_),.Y(_0098_));
NAND _1964_ (.A(_1385_),.B(_1513_),.Y(_1539_));
NAND _1965_ (.A(\mem[14] [12]),.B(_1514_),.Y(_1540_));
NAND _1966_ (.A(_1539_),.B(_1540_),.Y(_0099_));
NAND _1967_ (.A(_1388_),.B(_1513_),.Y(_1541_));
NAND _1968_ (.A(\mem[14] [13]),.B(_1514_),.Y(_1542_));
NAND _1969_ (.A(_1541_),.B(_1542_),.Y(_0100_));
NAND _1970_ (.A(_1391_),.B(_1513_),.Y(_1543_));
NAND _1971_ (.A(\mem[14] [14]),.B(_1514_),.Y(_1544_));
NAND _1972_ (.A(_1543_),.B(_1544_),.Y(_0101_));
NAND _1973_ (.A(_1393_),.B(_1513_),.Y(_1545_));
NAND _1974_ (.A(\mem[14] [15]),.B(_1514_),.Y(_1546_));
NAND _1975_ (.A(_1545_),.B(_1546_),.Y(_0102_));
NOR _1976_ (.A(_1399_),.B(_1442_),.Y(_1547_));
NAND _1977_ (.A(_1398_),.B(_1441_),.Y(_1548_));
NAND _1978_ (.A(_1402_),.B(_1547_),.Y(_1549_));
NAND _1979_ (.A(\mem[15] [0]),.B(_1548_),.Y(_1550_));
NAND _1980_ (.A(_1549_),.B(_1550_),.Y(_0112_));
NAND _1981_ (.A(_1405_),.B(_1547_),.Y(_1551_));
NAND _1982_ (.A(\mem[15] [1]),.B(_1548_),.Y(_1552_));
NAND _1983_ (.A(_1551_),.B(_1552_),.Y(_0119_));
NAND _1984_ (.A(_1408_),.B(_1547_),.Y(_1553_));
NAND _1985_ (.A(\mem[15] [2]),.B(_1548_),.Y(_1554_));
NAND _1986_ (.A(_1553_),.B(_1554_),.Y(_0120_));
NAND _1987_ (.A(_1357_),.B(_1547_),.Y(_1555_));
NAND _1988_ (.A(\mem[15] [3]),.B(_1548_),.Y(_1556_));
NAND _1989_ (.A(_1555_),.B(_1556_),.Y(_0121_));
NAND _1990_ (.A(_1361_),.B(_1547_),.Y(_1557_));
NAND _1991_ (.A(\mem[15] [4]),.B(_1548_),.Y(_1558_));
NAND _1992_ (.A(_1557_),.B(_1558_),.Y(_0122_));
NAND _1993_ (.A(_1364_),.B(_1547_),.Y(_1559_));
NAND _1994_ (.A(\mem[15] [5]),.B(_1548_),.Y(_1560_));
NAND _1995_ (.A(_1559_),.B(_1560_),.Y(_0123_));
NAND _1996_ (.A(_1367_),.B(_1547_),.Y(_1561_));
NAND _1997_ (.A(\mem[15] [6]),.B(_1548_),.Y(_1562_));
NAND _1998_ (.A(_1561_),.B(_1562_),.Y(_0124_));
NAND _1999_ (.A(_1370_),.B(_1547_),.Y(_1563_));
NAND _2000_ (.A(\mem[15] [7]),.B(_1548_),.Y(_1564_));
NAND _2001_ (.A(_1563_),.B(_1564_),.Y(_0125_));
NAND _2002_ (.A(_1372_),.B(_1547_),.Y(_1565_));
NAND _2003_ (.A(\mem[15] [8]),.B(_1548_),.Y(_1566_));
NAND _2004_ (.A(_1565_),.B(_1566_),.Y(_0126_));
NAND _2005_ (.A(_1375_),.B(_1547_),.Y(_1567_));
NAND _2006_ (.A(\mem[15] [9]),.B(_1548_),.Y(_1568_));
NAND _2007_ (.A(_1567_),.B(_1568_),.Y(_0127_));
NAND _2008_ (.A(_1379_),.B(_1547_),.Y(_1569_));
NAND _2009_ (.A(\mem[15] [10]),.B(_1548_),.Y(_1570_));
NAND _2010_ (.A(_1569_),.B(_1570_),.Y(_0113_));
NAND _2011_ (.A(_1382_),.B(_1547_),.Y(_1571_));
NAND _2012_ (.A(\mem[15] [11]),.B(_1548_),.Y(_1572_));
NAND _2013_ (.A(_1571_),.B(_1572_),.Y(_0114_));
NAND _2014_ (.A(_1385_),.B(_1547_),.Y(_1573_));
NAND _2015_ (.A(\mem[15] [12]),.B(_1548_),.Y(_1574_));
NAND _2016_ (.A(_1573_),.B(_1574_),.Y(_0115_));
NAND _2017_ (.A(_1388_),.B(_1547_),.Y(_1575_));
NAND _2018_ (.A(\mem[15] [13]),.B(_1548_),.Y(_1576_));
NAND _2019_ (.A(_1575_),.B(_1576_),.Y(_0116_));
NAND _2020_ (.A(_1391_),.B(_1547_),.Y(_1577_));
NAND _2021_ (.A(\mem[15] [14]),.B(_1548_),.Y(_1578_));
NAND _2022_ (.A(_1577_),.B(_1578_),.Y(_0117_));
NAND _2023_ (.A(_1393_),.B(_1547_),.Y(_1579_));
NAND _2024_ (.A(\mem[15] [15]),.B(_1548_),.Y(_1580_));
NAND _2025_ (.A(_1579_),.B(_1580_),.Y(_0118_));
NOR _2026_ (.A(_1279_),.B(_1331_),.Y(_1581_));
NAND _2027_ (.A(_1331_),.B(\mem[10] [0]),.Y(_1582_));
NAND _2028_ (.A(_1333_),.B(_1582_),.Y(_1583_));
NOR _2029_ (.A(_1581_),.B(_1583_),.Y(_1584_));
NOR _2030_ (.A(_1294_),.B(_1331_),.Y(_1585_));
NAND _2031_ (.A(\mem[11] [0]),.B(_1331_),.Y(_1586_));
NAND _2032_ (.A(read_addr[0]),.B(_1586_),.Y(_1587_));
NOR _2033_ (.A(_1585_),.B(_1587_),.Y(_1588_));
NOR _2034_ (.A(_1584_),.B(_1588_),.Y(_1589_));
NOR _2035_ (.A(_1332_),.B(_1589_),.Y(_1590_));
NOR _2036_ (.A(\mem[13] [0]),.B(_1331_),.Y(_1591_));
NOR _2037_ (.A(read_addr[2]),.B(\mem[9] [0]),.Y(_1592_));
NOR _2038_ (.A(_1591_),.B(_1592_),.Y(_1593_));
NOR _2039_ (.A(_1333_),.B(_1593_),.Y(_1594_));
NOR _2040_ (.A(\mem[12] [0]),.B(_1331_),.Y(_1595_));
NOR _2041_ (.A(read_addr[2]),.B(\mem[8] [0]),.Y(_1596_));
NOR _2042_ (.A(_1595_),.B(_1596_),.Y(_1597_));
NOR _2043_ (.A(read_addr[0]),.B(_1597_),.Y(_1598_));
NOR _2044_ (.A(_1594_),.B(_1598_),.Y(_1599_));
NOR _2045_ (.A(read_addr[1]),.B(_1599_),.Y(_1600_));
NOR _2046_ (.A(_1590_),.B(_1600_),.Y(_1601_));
NOR _2047_ (.A(_1330_),.B(_1601_),.Y(_1602_));
NAND _2048_ (.A(_1331_),.B(\mem[2] [0]),.Y(_1603_));
NAND _2049_ (.A(read_addr[2]),.B(\mem[6] [0]),.Y(_1604_));
NAND _2050_ (.A(_1603_),.B(_1604_),.Y(_1605_));
NOR _2051_ (.A(read_addr[0]),.B(_1605_),.Y(_1606_));
NOR _2052_ (.A(read_addr[2]),.B(_1334_),.Y(_1607_));
NAND _2053_ (.A(read_addr[2]),.B(\mem[7] [0]),.Y(_1608_));
NAND _2054_ (.A(read_addr[0]),.B(_1608_),.Y(_1609_));
NOR _2055_ (.A(_1607_),.B(_1609_),.Y(_1610_));
NOR _2056_ (.A(_1606_),.B(_1610_),.Y(_1611_));
NOR _2057_ (.A(_1332_),.B(_1611_),.Y(_1612_));
NOR _2058_ (.A(read_addr[2]),.B(\mem[1] [0]),.Y(_1613_));
NOR _2059_ (.A(_1331_),.B(\mem[5] [0]),.Y(_1614_));
NOR _2060_ (.A(_1613_),.B(_1614_),.Y(_1615_));
NOR _2061_ (.A(_1333_),.B(_1615_),.Y(_1616_));
NOR _2062_ (.A(read_addr[2]),.B(\mem[0] [0]),.Y(_1617_));
NOR _2063_ (.A(_1331_),.B(\mem[4] [0]),.Y(_1618_));
NOR _2064_ (.A(_1617_),.B(_1618_),.Y(_1619_));
NOR _2065_ (.A(read_addr[0]),.B(_1619_),.Y(_1620_));
NOR _2066_ (.A(_1616_),.B(_1620_),.Y(_1621_));
NOR _2067_ (.A(read_addr[1]),.B(_1621_),.Y(_1622_));
NOR _2068_ (.A(_1612_),.B(_1622_),.Y(_1623_));
NOR _2069_ (.A(read_addr[3]),.B(_1623_),.Y(_1624_));
NOR _2070_ (.A(_1602_),.B(_1624_),.Y(_0000_));
NOR _2071_ (.A(_1280_),.B(_1331_),.Y(_1625_));
NAND _2072_ (.A(_1331_),.B(\mem[10] [1]),.Y(_1626_));
NAND _2073_ (.A(_1333_),.B(_1626_),.Y(_1627_));
NOR _2074_ (.A(_1625_),.B(_1627_),.Y(_1628_));
NOR _2075_ (.A(_1295_),.B(_1331_),.Y(_1629_));
NAND _2076_ (.A(\mem[11] [1]),.B(_1331_),.Y(_1630_));
NAND _2077_ (.A(read_addr[0]),.B(_1630_),.Y(_0272_));
NOR _2078_ (.A(_1629_),.B(_0272_),.Y(_0273_));
NOR _2079_ (.A(_1628_),.B(_0273_),.Y(_0274_));
NOR _2080_ (.A(_1332_),.B(_0274_),.Y(_0275_));
NOR _2081_ (.A(read_addr[2]),.B(\mem[9] [1]),.Y(_0276_));
NOR _2082_ (.A(\mem[13] [1]),.B(_1331_),.Y(_0277_));
NOR _2083_ (.A(_0276_),.B(_0277_),.Y(_0278_));
NOR _2084_ (.A(_1333_),.B(_0278_),.Y(_0279_));
NOR _2085_ (.A(read_addr[2]),.B(\mem[8] [1]),.Y(_0280_));
NOR _2086_ (.A(\mem[12] [1]),.B(_1331_),.Y(_0281_));
NOR _2087_ (.A(_0280_),.B(_0281_),.Y(_0282_));
NOR _2088_ (.A(read_addr[0]),.B(_0282_),.Y(_0283_));
NOR _2089_ (.A(_0279_),.B(_0283_),.Y(_0284_));
NOR _2090_ (.A(read_addr[1]),.B(_0284_),.Y(_0285_));
NOR _2091_ (.A(_0275_),.B(_0285_),.Y(_0286_));
NOR _2092_ (.A(_1330_),.B(_0286_),.Y(_0287_));
NAND _2093_ (.A(_1331_),.B(\mem[2] [1]),.Y(_0288_));
NAND _2094_ (.A(read_addr[2]),.B(\mem[6] [1]),.Y(_0289_));
NAND _2095_ (.A(_0288_),.B(_0289_),.Y(_0290_));
NOR _2096_ (.A(read_addr[0]),.B(_0290_),.Y(_0291_));
NOR _2097_ (.A(read_addr[2]),.B(_1335_),.Y(_0292_));
NAND _2098_ (.A(read_addr[2]),.B(\mem[7] [1]),.Y(_0293_));
NAND _2099_ (.A(read_addr[0]),.B(_0293_),.Y(_0294_));
NOR _2100_ (.A(_0292_),.B(_0294_),.Y(_0295_));
NOR _2101_ (.A(_0291_),.B(_0295_),.Y(_0296_));
NOR _2102_ (.A(_1332_),.B(_0296_),.Y(_0297_));
NOR _2103_ (.A(read_addr[2]),.B(\mem[1] [1]),.Y(_0298_));
NOR _2104_ (.A(_1331_),.B(\mem[5] [1]),.Y(_0299_));
NOR _2105_ (.A(_0298_),.B(_0299_),.Y(_0300_));
NOR _2106_ (.A(_1333_),.B(_0300_),.Y(_0301_));
NOR _2107_ (.A(read_addr[2]),.B(\mem[0] [1]),.Y(_0302_));
NOR _2108_ (.A(_1331_),.B(\mem[4] [1]),.Y(_0303_));
NOR _2109_ (.A(_0302_),.B(_0303_),.Y(_0304_));
NOR _2110_ (.A(read_addr[0]),.B(_0304_),.Y(_0305_));
NOR _2111_ (.A(_0301_),.B(_0305_),.Y(_0306_));
NOR _2112_ (.A(read_addr[1]),.B(_0306_),.Y(_0307_));
NOR _2113_ (.A(_0297_),.B(_0307_),.Y(_0308_));
NOR _2114_ (.A(read_addr[3]),.B(_0308_),.Y(_0309_));
NOR _2115_ (.A(_0287_),.B(_0309_),.Y(_0007_));
NOR _2116_ (.A(_1331_),.B(\mem[7] [2]),.Y(_0310_));
NOR _2117_ (.A(read_addr[2]),.B(\mem[3] [2]),.Y(_0311_));
NOR _2118_ (.A(_0310_),.B(_0311_),.Y(_0312_));
NOR _2119_ (.A(_1333_),.B(_0312_),.Y(_0313_));
NOR _2120_ (.A(_1331_),.B(\mem[6] [2]),.Y(_0314_));
NOR _2121_ (.A(read_addr[2]),.B(\mem[2] [2]),.Y(_0315_));
NOR _2122_ (.A(_0314_),.B(_0315_),.Y(_0316_));
NOR _2123_ (.A(read_addr[0]),.B(_0316_),.Y(_0317_));
NOR _2124_ (.A(_0313_),.B(_0317_),.Y(_0318_));
NOR _2125_ (.A(_1332_),.B(_0318_),.Y(_0319_));
NOR _2126_ (.A(read_addr[2]),.B(\mem[1] [2]),.Y(_0320_));
NOR _2127_ (.A(_1331_),.B(\mem[5] [2]),.Y(_0321_));
NOR _2128_ (.A(_0320_),.B(_0321_),.Y(_0322_));
NOR _2129_ (.A(_1333_),.B(_0322_),.Y(_0323_));
NOR _2130_ (.A(read_addr[2]),.B(\mem[0] [2]),.Y(_0324_));
NOR _2131_ (.A(_1331_),.B(\mem[4] [2]),.Y(_0325_));
NOR _2132_ (.A(_0324_),.B(_0325_),.Y(_0326_));
NOR _2133_ (.A(read_addr[0]),.B(_0326_),.Y(_0327_));
NOR _2134_ (.A(_0323_),.B(_0327_),.Y(_0328_));
NOR _2135_ (.A(read_addr[1]),.B(_0328_),.Y(_0329_));
NOR _2136_ (.A(_0319_),.B(_0329_),.Y(_0330_));
NOR _2137_ (.A(read_addr[3]),.B(_0330_),.Y(_0331_));
NAND _2138_ (.A(\mem[12] [2]),.B(read_addr[2]),.Y(_0332_));
NAND _2139_ (.A(_1331_),.B(\mem[8] [2]),.Y(_0333_));
NAND _2140_ (.A(_0332_),.B(_0333_),.Y(_0334_));
NAND _2141_ (.A(_1333_),.B(_0334_),.Y(_0335_));
NAND _2142_ (.A(\mem[13] [2]),.B(read_addr[2]),.Y(_0336_));
NAND _2143_ (.A(_1331_),.B(\mem[9] [2]),.Y(_0337_));
NAND _2144_ (.A(_0336_),.B(_0337_),.Y(_0338_));
NAND _2145_ (.A(read_addr[0]),.B(_0338_),.Y(_0339_));
NAND _2146_ (.A(_0335_),.B(_0339_),.Y(_0340_));
NOR _2147_ (.A(read_addr[1]),.B(_0340_),.Y(_0341_));
NOR _2148_ (.A(\mem[15] [2]),.B(_1331_),.Y(_0342_));
NOR _2149_ (.A(\mem[11] [2]),.B(read_addr[2]),.Y(_0343_));
NOT _2150_ (.A(_0343_),.Y(_0344_));
NAND _2151_ (.A(read_addr[0]),.B(_0344_),.Y(_0345_));
NOR _2152_ (.A(_0342_),.B(_0345_),.Y(_0346_));
NAND _2153_ (.A(\mem[14] [2]),.B(read_addr[2]),.Y(_0347_));
NAND _2154_ (.A(_1331_),.B(\mem[10] [2]),.Y(_0348_));
NAND _2155_ (.A(_0347_),.B(_0348_),.Y(_0349_));
NAND _2156_ (.A(_1333_),.B(_0349_),.Y(_0350_));
NAND _2157_ (.A(read_addr[1]),.B(_0350_),.Y(_0351_));
NOR _2158_ (.A(_0346_),.B(_0351_),.Y(_0352_));
NOR _2159_ (.A(_0341_),.B(_0352_),.Y(_0353_));
NOR _2160_ (.A(_1330_),.B(_0353_),.Y(_0354_));
NOR _2161_ (.A(_0331_),.B(_0354_),.Y(_0008_));
NOR _2162_ (.A(_1281_),.B(_1331_),.Y(_0355_));
NAND _2163_ (.A(\mem[10] [3]),.B(_1331_),.Y(_0356_));
NAND _2164_ (.A(_1333_),.B(_0356_),.Y(_0357_));
NOR _2165_ (.A(_0355_),.B(_0357_),.Y(_0358_));
NOR _2166_ (.A(_1296_),.B(_1331_),.Y(_0359_));
NAND _2167_ (.A(\mem[11] [3]),.B(_1331_),.Y(_0360_));
NAND _2168_ (.A(read_addr[0]),.B(_0360_),.Y(_0361_));
NOR _2169_ (.A(_0359_),.B(_0361_),.Y(_0362_));
NOR _2170_ (.A(_0358_),.B(_0362_),.Y(_0363_));
NOR _2171_ (.A(_1330_),.B(_0363_),.Y(_0364_));
NOR _2172_ (.A(_1331_),.B(\mem[7] [3]),.Y(_0365_));
NOR _2173_ (.A(read_addr[2]),.B(\mem[3] [3]),.Y(_0366_));
NOR _2174_ (.A(_0365_),.B(_0366_),.Y(_0367_));
NOR _2175_ (.A(_1333_),.B(_0367_),.Y(_0368_));
NOR _2176_ (.A(_1331_),.B(\mem[6] [3]),.Y(_0369_));
NOR _2177_ (.A(read_addr[2]),.B(\mem[2] [3]),.Y(_0370_));
NOR _2178_ (.A(_0369_),.B(_0370_),.Y(_0371_));
NOR _2179_ (.A(read_addr[0]),.B(_0371_),.Y(_0372_));
NOR _2180_ (.A(_0368_),.B(_0372_),.Y(_0373_));
NOR _2181_ (.A(read_addr[3]),.B(_0373_),.Y(_0374_));
NOR _2182_ (.A(_0364_),.B(_0374_),.Y(_0375_));
NOR _2183_ (.A(_1332_),.B(_0375_),.Y(_0376_));
NOR _2184_ (.A(read_addr[2]),.B(_1339_),.Y(_0377_));
NAND _2185_ (.A(\mem[12] [3]),.B(read_addr[2]),.Y(_0378_));
NAND _2186_ (.A(_1333_),.B(_0378_),.Y(_0379_));
NOR _2187_ (.A(_0377_),.B(_0379_),.Y(_0380_));
NOR _2188_ (.A(read_addr[2]),.B(_1340_),.Y(_0381_));
NAND _2189_ (.A(\mem[13] [3]),.B(read_addr[2]),.Y(_0382_));
NAND _2190_ (.A(read_addr[0]),.B(_0382_),.Y(_0383_));
NOR _2191_ (.A(_0381_),.B(_0383_),.Y(_0384_));
NOR _2192_ (.A(_0380_),.B(_0384_),.Y(_0385_));
NOR _2193_ (.A(_1330_),.B(_0385_),.Y(_0386_));
NOR _2194_ (.A(read_addr[2]),.B(\mem[1] [3]),.Y(_0387_));
NOR _2195_ (.A(_1331_),.B(\mem[5] [3]),.Y(_0388_));
NOR _2196_ (.A(_0387_),.B(_0388_),.Y(_0389_));
NOR _2197_ (.A(_1333_),.B(_0389_),.Y(_0390_));
NOR _2198_ (.A(read_addr[2]),.B(\mem[0] [3]),.Y(_0391_));
NOR _2199_ (.A(_1331_),.B(\mem[4] [3]),.Y(_0392_));
NOR _2200_ (.A(_0391_),.B(_0392_),.Y(_0393_));
NOR _2201_ (.A(read_addr[0]),.B(_0393_),.Y(_0394_));
NOR _2202_ (.A(_0390_),.B(_0394_),.Y(_0395_));
NOR _2203_ (.A(read_addr[3]),.B(_0395_),.Y(_0396_));
NOR _2204_ (.A(_0386_),.B(_0396_),.Y(_0397_));
NOR _2205_ (.A(read_addr[1]),.B(_0397_),.Y(_0398_));
NOR _2206_ (.A(_0376_),.B(_0398_),.Y(_0009_));
NOR _2207_ (.A(_1282_),.B(_1331_),.Y(_0399_));
NAND _2208_ (.A(\mem[10] [4]),.B(_1331_),.Y(_0400_));
NAND _2209_ (.A(_1333_),.B(_0400_),.Y(_0401_));
NOR _2210_ (.A(_0399_),.B(_0401_),.Y(_0402_));
NOR _2211_ (.A(_1297_),.B(_1331_),.Y(_0403_));
NAND _2212_ (.A(\mem[11] [4]),.B(_1331_),.Y(_0404_));
NAND _2213_ (.A(read_addr[0]),.B(_0404_),.Y(_0405_));
NOR _2214_ (.A(_0403_),.B(_0405_),.Y(_0406_));
NOR _2215_ (.A(_0402_),.B(_0406_),.Y(_0407_));
NOR _2216_ (.A(_1330_),.B(_0407_),.Y(_0408_));
NOR _2217_ (.A(_1331_),.B(\mem[7] [4]),.Y(_0409_));
NOR _2218_ (.A(read_addr[2]),.B(\mem[3] [4]),.Y(_0410_));
NOR _2219_ (.A(_0409_),.B(_0410_),.Y(_0411_));
NOR _2220_ (.A(_1333_),.B(_0411_),.Y(_0412_));
NOR _2221_ (.A(_1331_),.B(\mem[6] [4]),.Y(_0413_));
NOR _2222_ (.A(read_addr[2]),.B(\mem[2] [4]),.Y(_0414_));
NOR _2223_ (.A(_0413_),.B(_0414_),.Y(_0415_));
NOR _2224_ (.A(read_addr[0]),.B(_0415_),.Y(_0416_));
NOR _2225_ (.A(_0412_),.B(_0416_),.Y(_0417_));
NOR _2226_ (.A(read_addr[3]),.B(_0417_),.Y(_0418_));
NOR _2227_ (.A(_0408_),.B(_0418_),.Y(_0419_));
NOR _2228_ (.A(_1332_),.B(_0419_),.Y(_0420_));
NAND _2229_ (.A(_1331_),.B(\mem[8] [4]),.Y(_0421_));
NAND _2230_ (.A(\mem[12] [4]),.B(read_addr[2]),.Y(_0422_));
NAND _2231_ (.A(_1331_),.B(\mem[9] [4]),.Y(_0423_));
NAND _2232_ (.A(\mem[13] [4]),.B(read_addr[2]),.Y(_0424_));
NAND _2233_ (.A(_0421_),.B(_0422_),.Y(_0425_));
NAND _2234_ (.A(_1333_),.B(_0425_),.Y(_0426_));
NAND _2235_ (.A(_0423_),.B(_0424_),.Y(_0427_));
NAND _2236_ (.A(read_addr[0]),.B(_0427_),.Y(_0428_));
NAND _2237_ (.A(_0426_),.B(_0428_),.Y(_0429_));
NOR _2238_ (.A(_1330_),.B(_0429_),.Y(_0430_));
NOR _2239_ (.A(read_addr[2]),.B(\mem[1] [4]),.Y(_0431_));
NOR _2240_ (.A(_1331_),.B(\mem[5] [4]),.Y(_0432_));
NOR _2241_ (.A(_0431_),.B(_0432_),.Y(_0433_));
NOR _2242_ (.A(_1333_),.B(_0433_),.Y(_0434_));
NOR _2243_ (.A(read_addr[2]),.B(\mem[0] [4]),.Y(_0435_));
NOR _2244_ (.A(_1331_),.B(\mem[4] [4]),.Y(_0436_));
NOR _2245_ (.A(_0435_),.B(_0436_),.Y(_0437_));
NOR _2246_ (.A(read_addr[0]),.B(_0437_),.Y(_0438_));
NOR _2247_ (.A(_0434_),.B(_0438_),.Y(_0439_));
NOR _2248_ (.A(read_addr[3]),.B(_0439_),.Y(_0440_));
NOR _2249_ (.A(_0430_),.B(_0440_),.Y(_0441_));
NOR _2250_ (.A(read_addr[1]),.B(_0441_),.Y(_0442_));
NOR _2251_ (.A(_0420_),.B(_0442_),.Y(_0010_));
NOR _2252_ (.A(_1283_),.B(_1331_),.Y(_0443_));
NAND _2253_ (.A(\mem[10] [5]),.B(_1331_),.Y(_0444_));
NAND _2254_ (.A(_1333_),.B(_0444_),.Y(_0445_));
NOR _2255_ (.A(_0443_),.B(_0445_),.Y(_0446_));
NOR _2256_ (.A(_1298_),.B(_1331_),.Y(_0447_));
NAND _2257_ (.A(\mem[11] [5]),.B(_1331_),.Y(_0448_));
NAND _2258_ (.A(read_addr[0]),.B(_0448_),.Y(_0449_));
NOR _2259_ (.A(_0447_),.B(_0449_),.Y(_0450_));
NOR _2260_ (.A(_0446_),.B(_0450_),.Y(_0451_));
NOR _2261_ (.A(_1330_),.B(_0451_),.Y(_0452_));
NOR _2262_ (.A(_1331_),.B(\mem[7] [5]),.Y(_0453_));
NOR _2263_ (.A(read_addr[2]),.B(\mem[3] [5]),.Y(_0454_));
NOR _2264_ (.A(_0453_),.B(_0454_),.Y(_0455_));
NOR _2265_ (.A(_1333_),.B(_0455_),.Y(_0456_));
NOR _2266_ (.A(_1331_),.B(\mem[6] [5]),.Y(_0457_));
NOR _2267_ (.A(read_addr[2]),.B(\mem[2] [5]),.Y(_0458_));
NOR _2268_ (.A(_0457_),.B(_0458_),.Y(_0459_));
NOR _2269_ (.A(read_addr[0]),.B(_0459_),.Y(_0460_));
NOR _2270_ (.A(_0456_),.B(_0460_),.Y(_0461_));
NOR _2271_ (.A(read_addr[3]),.B(_0461_),.Y(_0462_));
NOR _2272_ (.A(_0452_),.B(_0462_),.Y(_0463_));
NOR _2273_ (.A(_1332_),.B(_0463_),.Y(_0464_));
NOR _2274_ (.A(read_addr[2]),.B(_1341_),.Y(_0465_));
NAND _2275_ (.A(\mem[12] [5]),.B(read_addr[2]),.Y(_0466_));
NAND _2276_ (.A(_1333_),.B(_0466_),.Y(_0467_));
NOR _2277_ (.A(_0465_),.B(_0467_),.Y(_0468_));
NOR _2278_ (.A(read_addr[2]),.B(_1342_),.Y(_0469_));
NAND _2279_ (.A(\mem[13] [5]),.B(read_addr[2]),.Y(_0470_));
NAND _2280_ (.A(read_addr[0]),.B(_0470_),.Y(_0471_));
NOR _2281_ (.A(_0469_),.B(_0471_),.Y(_0472_));
NOR _2282_ (.A(_0468_),.B(_0472_),.Y(_0473_));
NOR _2283_ (.A(_1330_),.B(_0473_),.Y(_0474_));
NOR _2284_ (.A(read_addr[2]),.B(\mem[1] [5]),.Y(_0475_));
NOR _2285_ (.A(_1331_),.B(\mem[5] [5]),.Y(_0476_));
NOR _2286_ (.A(_0475_),.B(_0476_),.Y(_0477_));
NOR _2287_ (.A(_1333_),.B(_0477_),.Y(_0478_));
NOR _2288_ (.A(read_addr[2]),.B(\mem[0] [5]),.Y(_0479_));
NOR _2289_ (.A(_1331_),.B(\mem[4] [5]),.Y(_0480_));
NOR _2290_ (.A(_0479_),.B(_0480_),.Y(_0481_));
NOR _2291_ (.A(read_addr[0]),.B(_0481_),.Y(_0482_));
NOR _2292_ (.A(_0478_),.B(_0482_),.Y(_0483_));
NOR _2293_ (.A(read_addr[3]),.B(_0483_),.Y(_0484_));
NOR _2294_ (.A(_0474_),.B(_0484_),.Y(_0485_));
NOR _2295_ (.A(read_addr[1]),.B(_0485_),.Y(_0486_));
NOR _2296_ (.A(_0464_),.B(_0486_),.Y(_0011_));
NOR _2297_ (.A(_1284_),.B(_1331_),.Y(_0487_));
NAND _2298_ (.A(\mem[10] [6]),.B(_1331_),.Y(_0488_));
NAND _2299_ (.A(_1333_),.B(_0488_),.Y(_0489_));
NOR _2300_ (.A(_0487_),.B(_0489_),.Y(_0490_));
NOR _2301_ (.A(_1299_),.B(_1331_),.Y(_0491_));
NAND _2302_ (.A(\mem[11] [6]),.B(_1331_),.Y(_0492_));
NAND _2303_ (.A(read_addr[0]),.B(_0492_),.Y(_0493_));
NOR _2304_ (.A(_0491_),.B(_0493_),.Y(_0494_));
NOR _2305_ (.A(_0490_),.B(_0494_),.Y(_0495_));
NOR _2306_ (.A(_1330_),.B(_0495_),.Y(_0496_));
NOR _2307_ (.A(_1331_),.B(\mem[7] [6]),.Y(_0497_));
NOR _2308_ (.A(read_addr[2]),.B(\mem[3] [6]),.Y(_0498_));
NOR _2309_ (.A(_0497_),.B(_0498_),.Y(_0499_));
NOR _2310_ (.A(_1333_),.B(_0499_),.Y(_0500_));
NOR _2311_ (.A(_1331_),.B(\mem[6] [6]),.Y(_0501_));
NOR _2312_ (.A(read_addr[2]),.B(\mem[2] [6]),.Y(_0502_));
NOR _2313_ (.A(_0501_),.B(_0502_),.Y(_0503_));
NOR _2314_ (.A(read_addr[0]),.B(_0503_),.Y(_0504_));
NOR _2315_ (.A(_0500_),.B(_0504_),.Y(_0505_));
NOR _2316_ (.A(read_addr[3]),.B(_0505_),.Y(_0506_));
NOR _2317_ (.A(_0496_),.B(_0506_),.Y(_0507_));
NOR _2318_ (.A(_1332_),.B(_0507_),.Y(_0508_));
NAND _2319_ (.A(_1331_),.B(\mem[8] [6]),.Y(_0509_));
NAND _2320_ (.A(\mem[12] [6]),.B(read_addr[2]),.Y(_0510_));
NAND _2321_ (.A(_1331_),.B(\mem[9] [6]),.Y(_0511_));
NAND _2322_ (.A(\mem[13] [6]),.B(read_addr[2]),.Y(_0512_));
NAND _2323_ (.A(_0509_),.B(_0510_),.Y(_0513_));
NAND _2324_ (.A(_1333_),.B(_0513_),.Y(_0514_));
NAND _2325_ (.A(_0511_),.B(_0512_),.Y(_0515_));
NAND _2326_ (.A(read_addr[0]),.B(_0515_),.Y(_0516_));
NAND _2327_ (.A(_0514_),.B(_0516_),.Y(_0517_));
NOR _2328_ (.A(_1330_),.B(_0517_),.Y(_0518_));
NOR _2329_ (.A(read_addr[2]),.B(\mem[1] [6]),.Y(_0519_));
NOR _2330_ (.A(_1331_),.B(\mem[5] [6]),.Y(_0520_));
NOR _2331_ (.A(_0519_),.B(_0520_),.Y(_0521_));
NOR _2332_ (.A(_1333_),.B(_0521_),.Y(_0522_));
NOR _2333_ (.A(read_addr[2]),.B(\mem[0] [6]),.Y(_0523_));
NOR _2334_ (.A(_1331_),.B(\mem[4] [6]),.Y(_0524_));
NOR _2335_ (.A(_0523_),.B(_0524_),.Y(_0525_));
NOR _2336_ (.A(read_addr[0]),.B(_0525_),.Y(_0526_));
NOR _2337_ (.A(_0522_),.B(_0526_),.Y(_0527_));
NOR _2338_ (.A(read_addr[3]),.B(_0527_),.Y(_0528_));
NOR _2339_ (.A(_0518_),.B(_0528_),.Y(_0529_));
NOR _2340_ (.A(read_addr[1]),.B(_0529_),.Y(_0530_));
NOR _2341_ (.A(_0508_),.B(_0530_),.Y(_0012_));
NOR _2342_ (.A(_1285_),.B(_1331_),.Y(_0531_));
NAND _2343_ (.A(\mem[10] [7]),.B(_1331_),.Y(_0532_));
NAND _2344_ (.A(_1333_),.B(_0532_),.Y(_0533_));
NOR _2345_ (.A(_0531_),.B(_0533_),.Y(_0534_));
NOR _2346_ (.A(_1300_),.B(_1331_),.Y(_0535_));
NAND _2347_ (.A(\mem[11] [7]),.B(_1331_),.Y(_0536_));
NAND _2348_ (.A(read_addr[0]),.B(_0536_),.Y(_0537_));
NOR _2349_ (.A(_0535_),.B(_0537_),.Y(_0538_));
NOR _2350_ (.A(_0534_),.B(_0538_),.Y(_0539_));
NOR _2351_ (.A(_1330_),.B(_0539_),.Y(_0540_));
NOR _2352_ (.A(_1331_),.B(\mem[7] [7]),.Y(_0541_));
NOR _2353_ (.A(read_addr[2]),.B(\mem[3] [7]),.Y(_0542_));
NOR _2354_ (.A(_0541_),.B(_0542_),.Y(_0543_));
NOR _2355_ (.A(_1333_),.B(_0543_),.Y(_0544_));
NOR _2356_ (.A(_1331_),.B(\mem[6] [7]),.Y(_0545_));
NOR _2357_ (.A(read_addr[2]),.B(\mem[2] [7]),.Y(_0546_));
NOR _2358_ (.A(_0545_),.B(_0546_),.Y(_0547_));
NOR _2359_ (.A(read_addr[0]),.B(_0547_),.Y(_0548_));
NOR _2360_ (.A(_0544_),.B(_0548_),.Y(_0549_));
NOR _2361_ (.A(read_addr[3]),.B(_0549_),.Y(_0550_));
NOR _2362_ (.A(_0540_),.B(_0550_),.Y(_0551_));
NOR _2363_ (.A(_1332_),.B(_0551_),.Y(_0552_));
NOR _2364_ (.A(read_addr[2]),.B(_1343_),.Y(_0553_));
NAND _2365_ (.A(\mem[12] [7]),.B(read_addr[2]),.Y(_0554_));
NAND _2366_ (.A(_1333_),.B(_0554_),.Y(_0555_));
NOR _2367_ (.A(_0553_),.B(_0555_),.Y(_0556_));
NOR _2368_ (.A(read_addr[2]),.B(_1344_),.Y(_0557_));
NAND _2369_ (.A(\mem[13] [7]),.B(read_addr[2]),.Y(_0558_));
NAND _2370_ (.A(read_addr[0]),.B(_0558_),.Y(_0559_));
NOR _2371_ (.A(_0557_),.B(_0559_),.Y(_0560_));
NOR _2372_ (.A(_0556_),.B(_0560_),.Y(_0561_));
NOR _2373_ (.A(_1330_),.B(_0561_),.Y(_0562_));
NOR _2374_ (.A(read_addr[2]),.B(\mem[1] [7]),.Y(_0563_));
NOR _2375_ (.A(_1331_),.B(\mem[5] [7]),.Y(_0564_));
NOR _2376_ (.A(_0563_),.B(_0564_),.Y(_0565_));
NOR _2377_ (.A(_1333_),.B(_0565_),.Y(_0566_));
NOR _2378_ (.A(read_addr[2]),.B(\mem[0] [7]),.Y(_0567_));
NOR _2379_ (.A(_1331_),.B(\mem[4] [7]),.Y(_0568_));
NOR _2380_ (.A(_0567_),.B(_0568_),.Y(_0569_));
NOR _2381_ (.A(read_addr[0]),.B(_0569_),.Y(_0570_));
NOR _2382_ (.A(_0566_),.B(_0570_),.Y(_0571_));
NOR _2383_ (.A(read_addr[3]),.B(_0571_),.Y(_0572_));
NOR _2384_ (.A(_0562_),.B(_0572_),.Y(_0573_));
NOR _2385_ (.A(read_addr[1]),.B(_0573_),.Y(_0574_));
NOR _2386_ (.A(_0552_),.B(_0574_),.Y(_0013_));
NOR _2387_ (.A(_1286_),.B(_1331_),.Y(_0575_));
NAND _2388_ (.A(\mem[10] [8]),.B(_1331_),.Y(_0576_));
NAND _2389_ (.A(_1333_),.B(_0576_),.Y(_0577_));
NOR _2390_ (.A(_0575_),.B(_0577_),.Y(_0578_));
NOR _2391_ (.A(_1301_),.B(_1331_),.Y(_0579_));
NAND _2392_ (.A(\mem[11] [8]),.B(_1331_),.Y(_0580_));
NAND _2393_ (.A(read_addr[0]),.B(_0580_),.Y(_0581_));
NOR _2394_ (.A(_0579_),.B(_0581_),.Y(_0582_));
NOR _2395_ (.A(_0578_),.B(_0582_),.Y(_0583_));
NOR _2396_ (.A(_1330_),.B(_0583_),.Y(_0584_));
NOR _2397_ (.A(_1331_),.B(\mem[7] [8]),.Y(_0585_));
NOR _2398_ (.A(read_addr[2]),.B(\mem[3] [8]),.Y(_0586_));
NOR _2399_ (.A(_0585_),.B(_0586_),.Y(_0587_));
NOR _2400_ (.A(_1333_),.B(_0587_),.Y(_0588_));
NOR _2401_ (.A(_1331_),.B(\mem[6] [8]),.Y(_0589_));
NOR _2402_ (.A(read_addr[2]),.B(\mem[2] [8]),.Y(_0590_));
NOR _2403_ (.A(_0589_),.B(_0590_),.Y(_0591_));
NOR _2404_ (.A(read_addr[0]),.B(_0591_),.Y(_0592_));
NOR _2405_ (.A(_0588_),.B(_0592_),.Y(_0593_));
NOR _2406_ (.A(read_addr[3]),.B(_0593_),.Y(_0594_));
NOR _2407_ (.A(_0584_),.B(_0594_),.Y(_0595_));
NOR _2408_ (.A(_1332_),.B(_0595_),.Y(_0596_));
NAND _2409_ (.A(_1331_),.B(\mem[8] [8]),.Y(_0597_));
NAND _2410_ (.A(\mem[12] [8]),.B(read_addr[2]),.Y(_0598_));
NAND _2411_ (.A(_1331_),.B(\mem[9] [8]),.Y(_0599_));
NAND _2412_ (.A(\mem[13] [8]),.B(read_addr[2]),.Y(_0600_));
NAND _2413_ (.A(_0597_),.B(_0598_),.Y(_0601_));
NAND _2414_ (.A(_1333_),.B(_0601_),.Y(_0602_));
NAND _2415_ (.A(_0599_),.B(_0600_),.Y(_0603_));
NAND _2416_ (.A(read_addr[0]),.B(_0603_),.Y(_0604_));
NAND _2417_ (.A(_0602_),.B(_0604_),.Y(_0605_));
NOR _2418_ (.A(_1330_),.B(_0605_),.Y(_0606_));
NOR _2419_ (.A(read_addr[2]),.B(\mem[1] [8]),.Y(_0607_));
NOR _2420_ (.A(_1331_),.B(\mem[5] [8]),.Y(_0608_));
NOR _2421_ (.A(_0607_),.B(_0608_),.Y(_0609_));
NOR _2422_ (.A(_1333_),.B(_0609_),.Y(_0610_));
NOR _2423_ (.A(read_addr[2]),.B(\mem[0] [8]),.Y(_0611_));
NOR _2424_ (.A(_1331_),.B(\mem[4] [8]),.Y(_0612_));
NOR _2425_ (.A(_0611_),.B(_0612_),.Y(_0613_));
NOR _2426_ (.A(read_addr[0]),.B(_0613_),.Y(_0614_));
NOR _2427_ (.A(_0610_),.B(_0614_),.Y(_0615_));
NOR _2428_ (.A(read_addr[3]),.B(_0615_),.Y(_0616_));
NOR _2429_ (.A(_0606_),.B(_0616_),.Y(_0617_));
NOR _2430_ (.A(read_addr[1]),.B(_0617_),.Y(_0618_));
NOR _2431_ (.A(_0596_),.B(_0618_),.Y(_0014_));
NOR _2432_ (.A(_1287_),.B(_1331_),.Y(_0619_));
NAND _2433_ (.A(\mem[10] [9]),.B(_1331_),.Y(_0620_));
NAND _2434_ (.A(_1333_),.B(_0620_),.Y(_0621_));
NOR _2435_ (.A(_0619_),.B(_0621_),.Y(_0622_));
NOR _2436_ (.A(_1302_),.B(_1331_),.Y(_0623_));
NAND _2437_ (.A(\mem[11] [9]),.B(_1331_),.Y(_0624_));
NAND _2438_ (.A(read_addr[0]),.B(_0624_),.Y(_0625_));
NOR _2439_ (.A(_0623_),.B(_0625_),.Y(_0626_));
NOR _2440_ (.A(_0622_),.B(_0626_),.Y(_0627_));
NOR _2441_ (.A(_1332_),.B(_0627_),.Y(_0628_));
NOR _2442_ (.A(read_addr[2]),.B(\mem[9] [9]),.Y(_0629_));
NOR _2443_ (.A(\mem[13] [9]),.B(_1331_),.Y(_0630_));
NOR _2444_ (.A(_0629_),.B(_0630_),.Y(_0631_));
NOR _2445_ (.A(_1333_),.B(_0631_),.Y(_0632_));
NOR _2446_ (.A(read_addr[2]),.B(\mem[8] [9]),.Y(_0633_));
NOR _2447_ (.A(\mem[12] [9]),.B(_1331_),.Y(_0634_));
NOR _2448_ (.A(_0633_),.B(_0634_),.Y(_0635_));
NOR _2449_ (.A(read_addr[0]),.B(_0635_),.Y(_0636_));
NOR _2450_ (.A(_0632_),.B(_0636_),.Y(_0637_));
NOR _2451_ (.A(read_addr[1]),.B(_0637_),.Y(_0638_));
NOR _2452_ (.A(_0628_),.B(_0638_),.Y(_0639_));
NOR _2453_ (.A(_1330_),.B(_0639_),.Y(_0640_));
NAND _2454_ (.A(_1331_),.B(\mem[2] [9]),.Y(_0641_));
NAND _2455_ (.A(read_addr[2]),.B(\mem[6] [9]),.Y(_0642_));
NAND _2456_ (.A(_0641_),.B(_0642_),.Y(_0643_));
NOR _2457_ (.A(read_addr[0]),.B(_0643_),.Y(_0644_));
NOR _2458_ (.A(read_addr[2]),.B(_1336_),.Y(_0645_));
NAND _2459_ (.A(read_addr[2]),.B(\mem[7] [9]),.Y(_0646_));
NAND _2460_ (.A(read_addr[0]),.B(_0646_),.Y(_0647_));
NOR _2461_ (.A(_0645_),.B(_0647_),.Y(_0648_));
NOR _2462_ (.A(_0644_),.B(_0648_),.Y(_0649_));
NOR _2463_ (.A(_1332_),.B(_0649_),.Y(_0650_));
NOR _2464_ (.A(read_addr[2]),.B(\mem[1] [9]),.Y(_0651_));
NOR _2465_ (.A(_1331_),.B(\mem[5] [9]),.Y(_0652_));
NOR _2466_ (.A(_0651_),.B(_0652_),.Y(_0653_));
NOR _2467_ (.A(_1333_),.B(_0653_),.Y(_0654_));
NOR _2468_ (.A(read_addr[2]),.B(\mem[0] [9]),.Y(_0655_));
NOR _2469_ (.A(_1331_),.B(\mem[4] [9]),.Y(_0656_));
NOR _2470_ (.A(_0655_),.B(_0656_),.Y(_0657_));
NOR _2471_ (.A(read_addr[0]),.B(_0657_),.Y(_0658_));
NOR _2472_ (.A(_0654_),.B(_0658_),.Y(_0659_));
NOR _2473_ (.A(read_addr[1]),.B(_0659_),.Y(_0660_));
NOR _2474_ (.A(_0650_),.B(_0660_),.Y(_0661_));
NOR _2475_ (.A(read_addr[3]),.B(_0661_),.Y(_0662_));
NOR _2476_ (.A(_0640_),.B(_0662_),.Y(_0015_));
NOR _2477_ (.A(_1288_),.B(_1331_),.Y(_0663_));
NAND _2478_ (.A(\mem[10] [10]),.B(_1331_),.Y(_0664_));
NAND _2479_ (.A(_1333_),.B(_0664_),.Y(_0665_));
NOR _2480_ (.A(_0663_),.B(_0665_),.Y(_0666_));
NOR _2481_ (.A(_1303_),.B(_1331_),.Y(_0667_));
NAND _2482_ (.A(\mem[11] [10]),.B(_1331_),.Y(_0668_));
NAND _2483_ (.A(read_addr[0]),.B(_0668_),.Y(_0669_));
NOR _2484_ (.A(_0667_),.B(_0669_),.Y(_0670_));
NOR _2485_ (.A(_0666_),.B(_0670_),.Y(_0671_));
NOR _2486_ (.A(_1332_),.B(_0671_),.Y(_0672_));
NOR _2487_ (.A(read_addr[2]),.B(\mem[9] [10]),.Y(_0673_));
NOR _2488_ (.A(\mem[13] [10]),.B(_1331_),.Y(_0674_));
NOR _2489_ (.A(_0673_),.B(_0674_),.Y(_0675_));
NOR _2490_ (.A(_1333_),.B(_0675_),.Y(_0676_));
NOR _2491_ (.A(read_addr[2]),.B(\mem[8] [10]),.Y(_0677_));
NOR _2492_ (.A(\mem[12] [10]),.B(_1331_),.Y(_0678_));
NOR _2493_ (.A(_0677_),.B(_0678_),.Y(_0679_));
NOR _2494_ (.A(read_addr[0]),.B(_0679_),.Y(_0680_));
NOR _2495_ (.A(_0676_),.B(_0680_),.Y(_0681_));
NOR _2496_ (.A(read_addr[1]),.B(_0681_),.Y(_0682_));
NOR _2497_ (.A(_0672_),.B(_0682_),.Y(_0683_));
NOR _2498_ (.A(_1330_),.B(_0683_),.Y(_0684_));
NAND _2499_ (.A(_1331_),.B(\mem[2] [10]),.Y(_0685_));
NAND _2500_ (.A(read_addr[2]),.B(\mem[6] [10]),.Y(_0686_));
NAND _2501_ (.A(_0685_),.B(_0686_),.Y(_0687_));
NOR _2502_ (.A(read_addr[0]),.B(_0687_),.Y(_0688_));
NOR _2503_ (.A(read_addr[2]),.B(_1337_),.Y(_0689_));
NAND _2504_ (.A(read_addr[2]),.B(\mem[7] [10]),.Y(_0690_));
NAND _2505_ (.A(read_addr[0]),.B(_0690_),.Y(_0691_));
NOR _2506_ (.A(_0689_),.B(_0691_),.Y(_0692_));
NOR _2507_ (.A(_0688_),.B(_0692_),.Y(_0693_));
NOR _2508_ (.A(_1332_),.B(_0693_),.Y(_0694_));
NOR _2509_ (.A(read_addr[2]),.B(\mem[1] [10]),.Y(_0695_));
NOR _2510_ (.A(_1331_),.B(\mem[5] [10]),.Y(_0696_));
NOR _2511_ (.A(_0695_),.B(_0696_),.Y(_0697_));
NOR _2512_ (.A(_1333_),.B(_0697_),.Y(_0698_));
NOR _2513_ (.A(read_addr[2]),.B(\mem[0] [10]),.Y(_0699_));
NOR _2514_ (.A(_1331_),.B(\mem[4] [10]),.Y(_0700_));
NOR _2515_ (.A(_0699_),.B(_0700_),.Y(_0701_));
NOR _2516_ (.A(read_addr[0]),.B(_0701_),.Y(_0702_));
NOR _2517_ (.A(_0698_),.B(_0702_),.Y(_0703_));
NOR _2518_ (.A(read_addr[1]),.B(_0703_),.Y(_0704_));
NOR _2519_ (.A(_0694_),.B(_0704_),.Y(_0705_));
NOR _2520_ (.A(read_addr[3]),.B(_0705_),.Y(_0706_));
NOR _2521_ (.A(_0684_),.B(_0706_),.Y(_0001_));
NOR _2522_ (.A(_1289_),.B(_1331_),.Y(_0707_));
NAND _2523_ (.A(\mem[10] [11]),.B(_1331_),.Y(_0708_));
NAND _2524_ (.A(_1333_),.B(_0708_),.Y(_0709_));
NOR _2525_ (.A(_0707_),.B(_0709_),.Y(_0710_));
NOR _2526_ (.A(_1304_),.B(_1331_),.Y(_0711_));
NAND _2527_ (.A(\mem[11] [11]),.B(_1331_),.Y(_0712_));
NAND _2528_ (.A(read_addr[0]),.B(_0712_),.Y(_0713_));
NOR _2529_ (.A(_0711_),.B(_0713_),.Y(_0714_));
NOR _2530_ (.A(_0710_),.B(_0714_),.Y(_0715_));
NOR _2531_ (.A(_1330_),.B(_0715_),.Y(_0716_));
NOR _2532_ (.A(_1331_),.B(\mem[7] [11]),.Y(_0717_));
NOR _2533_ (.A(read_addr[2]),.B(\mem[3] [11]),.Y(_0718_));
NOR _2534_ (.A(_0717_),.B(_0718_),.Y(_0719_));
NOR _2535_ (.A(_1333_),.B(_0719_),.Y(_0720_));
NOR _2536_ (.A(_1331_),.B(\mem[6] [11]),.Y(_0721_));
NOR _2537_ (.A(read_addr[2]),.B(\mem[2] [11]),.Y(_0722_));
NOR _2538_ (.A(_0721_),.B(_0722_),.Y(_0723_));
NOR _2539_ (.A(read_addr[0]),.B(_0723_),.Y(_0724_));
NOR _2540_ (.A(_0720_),.B(_0724_),.Y(_0725_));
NOR _2541_ (.A(read_addr[3]),.B(_0725_),.Y(_0726_));
NOR _2542_ (.A(_0716_),.B(_0726_),.Y(_0727_));
NOR _2543_ (.A(_1332_),.B(_0727_),.Y(_0728_));
NAND _2544_ (.A(_1331_),.B(\mem[8] [11]),.Y(_0729_));
NAND _2545_ (.A(\mem[12] [11]),.B(read_addr[2]),.Y(_0730_));
NAND _2546_ (.A(_1331_),.B(\mem[9] [11]),.Y(_0731_));
NAND _2547_ (.A(\mem[13] [11]),.B(read_addr[2]),.Y(_0732_));
NAND _2548_ (.A(_0729_),.B(_0730_),.Y(_0733_));
NAND _2549_ (.A(_1333_),.B(_0733_),.Y(_0734_));
NAND _2550_ (.A(_0731_),.B(_0732_),.Y(_0735_));
NAND _2551_ (.A(read_addr[0]),.B(_0735_),.Y(_0736_));
NAND _2552_ (.A(_0734_),.B(_0736_),.Y(_0737_));
NOR _2553_ (.A(_1330_),.B(_0737_),.Y(_0738_));
NOR _2554_ (.A(read_addr[2]),.B(\mem[1] [11]),.Y(_0739_));
NOR _2555_ (.A(_1331_),.B(\mem[5] [11]),.Y(_0740_));
NOR _2556_ (.A(_0739_),.B(_0740_),.Y(_0741_));
NOR _2557_ (.A(_1333_),.B(_0741_),.Y(_0742_));
NOR _2558_ (.A(read_addr[2]),.B(\mem[0] [11]),.Y(_0743_));
NOR _2559_ (.A(_1331_),.B(\mem[4] [11]),.Y(_0744_));
NOR _2560_ (.A(_0743_),.B(_0744_),.Y(_0745_));
NOR _2561_ (.A(read_addr[0]),.B(_0745_),.Y(_0746_));
NOR _2562_ (.A(_0742_),.B(_0746_),.Y(_0747_));
NOR _2563_ (.A(read_addr[3]),.B(_0747_),.Y(_0748_));
NOR _2564_ (.A(_0738_),.B(_0748_),.Y(_0749_));
NOR _2565_ (.A(read_addr[1]),.B(_0749_),.Y(_0750_));
NOR _2566_ (.A(_0728_),.B(_0750_),.Y(_0002_));
NOR _2567_ (.A(_1290_),.B(_1331_),.Y(_0751_));
NAND _2568_ (.A(\mem[10] [12]),.B(_1331_),.Y(_0752_));
NAND _2569_ (.A(_1333_),.B(_0752_),.Y(_0753_));
NOR _2570_ (.A(_0751_),.B(_0753_),.Y(_0754_));
NOR _2571_ (.A(_1305_),.B(_1331_),.Y(_0755_));
NAND _2572_ (.A(\mem[11] [12]),.B(_1331_),.Y(_0756_));
NAND _2573_ (.A(read_addr[0]),.B(_0756_),.Y(_0757_));
NOR _2574_ (.A(_0755_),.B(_0757_),.Y(_0758_));
NOR _2575_ (.A(_0754_),.B(_0758_),.Y(_0759_));
NOR _2576_ (.A(_1330_),.B(_0759_),.Y(_0760_));
NOR _2577_ (.A(_1331_),.B(\mem[7] [12]),.Y(_0761_));
NOR _2578_ (.A(read_addr[2]),.B(\mem[3] [12]),.Y(_0762_));
NOR _2579_ (.A(_0761_),.B(_0762_),.Y(_0763_));
NOR _2580_ (.A(_1333_),.B(_0763_),.Y(_0764_));
NOR _2581_ (.A(_1331_),.B(\mem[6] [12]),.Y(_0765_));
NOR _2582_ (.A(read_addr[2]),.B(\mem[2] [12]),.Y(_0766_));
NOR _2583_ (.A(_0765_),.B(_0766_),.Y(_0767_));
NOR _2584_ (.A(read_addr[0]),.B(_0767_),.Y(_0768_));
NOR _2585_ (.A(_0764_),.B(_0768_),.Y(_0769_));
NOR _2586_ (.A(read_addr[3]),.B(_0769_),.Y(_0770_));
NOR _2587_ (.A(_0760_),.B(_0770_),.Y(_0771_));
NOR _2588_ (.A(_1332_),.B(_0771_),.Y(_0772_));
NAND _2589_ (.A(_1331_),.B(\mem[8] [12]),.Y(_0773_));
NAND _2590_ (.A(\mem[12] [12]),.B(read_addr[2]),.Y(_0774_));
NAND _2591_ (.A(_1331_),.B(\mem[9] [12]),.Y(_0775_));
NAND _2592_ (.A(\mem[13] [12]),.B(read_addr[2]),.Y(_0776_));
NAND _2593_ (.A(_0773_),.B(_0774_),.Y(_0777_));
NAND _2594_ (.A(_1333_),.B(_0777_),.Y(_0778_));
NAND _2595_ (.A(_0775_),.B(_0776_),.Y(_0779_));
NAND _2596_ (.A(read_addr[0]),.B(_0779_),.Y(_0780_));
NAND _2597_ (.A(_0778_),.B(_0780_),.Y(_0781_));
NOR _2598_ (.A(_1330_),.B(_0781_),.Y(_0782_));
NOR _2599_ (.A(read_addr[2]),.B(\mem[1] [12]),.Y(_0783_));
NOR _2600_ (.A(_1331_),.B(\mem[5] [12]),.Y(_0784_));
NOR _2601_ (.A(_0783_),.B(_0784_),.Y(_0785_));
NOR _2602_ (.A(_1333_),.B(_0785_),.Y(_0786_));
NOR _2603_ (.A(read_addr[2]),.B(\mem[0] [12]),.Y(_0787_));
NOR _2604_ (.A(_1331_),.B(\mem[4] [12]),.Y(_0788_));
NOR _2605_ (.A(_0787_),.B(_0788_),.Y(_0789_));
NOR _2606_ (.A(read_addr[0]),.B(_0789_),.Y(_0790_));
NOR _2607_ (.A(_0786_),.B(_0790_),.Y(_0791_));
NOR _2608_ (.A(read_addr[3]),.B(_0791_),.Y(_0792_));
NOR _2609_ (.A(_0782_),.B(_0792_),.Y(_0793_));
NOR _2610_ (.A(read_addr[1]),.B(_0793_),.Y(_0794_));
NOR _2611_ (.A(_0772_),.B(_0794_),.Y(_0003_));
NOR _2612_ (.A(_1291_),.B(_1331_),.Y(_0795_));
NAND _2613_ (.A(\mem[10] [13]),.B(_1331_),.Y(_0796_));
NAND _2614_ (.A(_1333_),.B(_0796_),.Y(_0797_));
NOR _2615_ (.A(_0795_),.B(_0797_),.Y(_0798_));
NOR _2616_ (.A(_1306_),.B(_1331_),.Y(_0799_));
NAND _2617_ (.A(\mem[11] [13]),.B(_1331_),.Y(_0800_));
NAND _2618_ (.A(read_addr[0]),.B(_0800_),.Y(_0801_));
NOR _2619_ (.A(_0799_),.B(_0801_),.Y(_0802_));
NOR _2620_ (.A(_0798_),.B(_0802_),.Y(_0803_));
NOR _2621_ (.A(_1330_),.B(_0803_),.Y(_0804_));
NOR _2622_ (.A(_1331_),.B(\mem[7] [13]),.Y(_0805_));
NOR _2623_ (.A(read_addr[2]),.B(\mem[3] [13]),.Y(_0806_));
NOR _2624_ (.A(_0805_),.B(_0806_),.Y(_0807_));
NOR _2625_ (.A(_1333_),.B(_0807_),.Y(_0808_));
NOR _2626_ (.A(_1331_),.B(\mem[6] [13]),.Y(_0809_));
NOR _2627_ (.A(read_addr[2]),.B(\mem[2] [13]),.Y(_0810_));
NOR _2628_ (.A(_0809_),.B(_0810_),.Y(_0811_));
NOR _2629_ (.A(read_addr[0]),.B(_0811_),.Y(_0812_));
NOR _2630_ (.A(_0808_),.B(_0812_),.Y(_0813_));
NOR _2631_ (.A(read_addr[3]),.B(_0813_),.Y(_0814_));
NOR _2632_ (.A(_0804_),.B(_0814_),.Y(_0815_));
NOR _2633_ (.A(_1332_),.B(_0815_),.Y(_0816_));
NAND _2634_ (.A(_1331_),.B(\mem[8] [13]),.Y(_0817_));
NAND _2635_ (.A(\mem[12] [13]),.B(read_addr[2]),.Y(_0818_));
NAND _2636_ (.A(_1331_),.B(\mem[9] [13]),.Y(_0819_));
NAND _2637_ (.A(\mem[13] [13]),.B(read_addr[2]),.Y(_0820_));
NAND _2638_ (.A(_0817_),.B(_0818_),.Y(_0821_));
NAND _2639_ (.A(_1333_),.B(_0821_),.Y(_0822_));
NAND _2640_ (.A(_0819_),.B(_0820_),.Y(_0823_));
NAND _2641_ (.A(read_addr[0]),.B(_0823_),.Y(_0824_));
NAND _2642_ (.A(_0822_),.B(_0824_),.Y(_0825_));
NOR _2643_ (.A(_1330_),.B(_0825_),.Y(_0826_));
NOR _2644_ (.A(read_addr[2]),.B(\mem[1] [13]),.Y(_0827_));
NOR _2645_ (.A(_1331_),.B(\mem[5] [13]),.Y(_0828_));
NOR _2646_ (.A(_0827_),.B(_0828_),.Y(_0829_));
NOR _2647_ (.A(_1333_),.B(_0829_),.Y(_0830_));
NOR _2648_ (.A(read_addr[2]),.B(\mem[0] [13]),.Y(_0831_));
NOR _2649_ (.A(_1331_),.B(\mem[4] [13]),.Y(_0832_));
NOR _2650_ (.A(_0831_),.B(_0832_),.Y(_0833_));
NOR _2651_ (.A(read_addr[0]),.B(_0833_),.Y(_0834_));
NOR _2652_ (.A(_0830_),.B(_0834_),.Y(_0835_));
NOR _2653_ (.A(read_addr[3]),.B(_0835_),.Y(_0836_));
NOR _2654_ (.A(_0826_),.B(_0836_),.Y(_0837_));
NOR _2655_ (.A(read_addr[1]),.B(_0837_),.Y(_0838_));
NOR _2656_ (.A(_0816_),.B(_0838_),.Y(_0004_));
NOR _2657_ (.A(_1292_),.B(_1331_),.Y(_0839_));
NAND _2658_ (.A(\mem[10] [14]),.B(_1331_),.Y(_0840_));
NAND _2659_ (.A(_1333_),.B(_0840_),.Y(_0841_));
NOR _2660_ (.A(_0839_),.B(_0841_),.Y(_0842_));
NOR _2661_ (.A(_1307_),.B(_1331_),.Y(_0843_));
NAND _2662_ (.A(\mem[11] [14]),.B(_1331_),.Y(_0844_));
NAND _2663_ (.A(read_addr[0]),.B(_0844_),.Y(_0845_));
NOR _2664_ (.A(_0843_),.B(_0845_),.Y(_0846_));
NOR _2665_ (.A(_0842_),.B(_0846_),.Y(_0847_));
NOR _2666_ (.A(_1332_),.B(_0847_),.Y(_0848_));
NOR _2667_ (.A(\mem[13] [14]),.B(_1331_),.Y(_0849_));
NOR _2668_ (.A(read_addr[2]),.B(\mem[9] [14]),.Y(_0850_));
NOR _2669_ (.A(_0849_),.B(_0850_),.Y(_0851_));
NOR _2670_ (.A(_1333_),.B(_0851_),.Y(_0852_));
NOR _2671_ (.A(\mem[12] [14]),.B(_1331_),.Y(_0853_));
NOR _2672_ (.A(read_addr[2]),.B(\mem[8] [14]),.Y(_0854_));
NOR _2673_ (.A(_0853_),.B(_0854_),.Y(_0855_));
NOR _2674_ (.A(read_addr[0]),.B(_0855_),.Y(_0856_));
NOR _2675_ (.A(_0852_),.B(_0856_),.Y(_0857_));
NOR _2676_ (.A(read_addr[1]),.B(_0857_),.Y(_0858_));
NOR _2677_ (.A(_0848_),.B(_0858_),.Y(_0859_));
NOR _2678_ (.A(_1330_),.B(_0859_),.Y(_0860_));
NAND _2679_ (.A(_1331_),.B(\mem[2] [14]),.Y(_0861_));
NAND _2680_ (.A(read_addr[2]),.B(\mem[6] [14]),.Y(_0862_));
NAND _2681_ (.A(_0861_),.B(_0862_),.Y(_0863_));
NOR _2682_ (.A(read_addr[0]),.B(_0863_),.Y(_0864_));
NOR _2683_ (.A(read_addr[2]),.B(_1338_),.Y(_0865_));
NAND _2684_ (.A(read_addr[2]),.B(\mem[7] [14]),.Y(_0866_));
NAND _2685_ (.A(read_addr[0]),.B(_0866_),.Y(_0867_));
NOR _2686_ (.A(_0865_),.B(_0867_),.Y(_0868_));
NOR _2687_ (.A(_0864_),.B(_0868_),.Y(_0869_));
NOR _2688_ (.A(_1332_),.B(_0869_),.Y(_0870_));
NOR _2689_ (.A(read_addr[2]),.B(\mem[1] [14]),.Y(_0871_));
NOR _2690_ (.A(_1331_),.B(\mem[5] [14]),.Y(_0872_));
NOR _2691_ (.A(_0871_),.B(_0872_),.Y(_0873_));
NOR _2692_ (.A(_1333_),.B(_0873_),.Y(_0874_));
NOR _2693_ (.A(read_addr[2]),.B(\mem[0] [14]),.Y(_0875_));
NOR _2694_ (.A(_1331_),.B(\mem[4] [14]),.Y(_0876_));
NOR _2695_ (.A(_0875_),.B(_0876_),.Y(_0877_));
NOR _2696_ (.A(read_addr[0]),.B(_0877_),.Y(_0878_));
NOR _2697_ (.A(_0874_),.B(_0878_),.Y(_0879_));
NOR _2698_ (.A(read_addr[1]),.B(_0879_),.Y(_0880_));
NOR _2699_ (.A(_0870_),.B(_0880_),.Y(_0881_));
NOR _2700_ (.A(read_addr[3]),.B(_0881_),.Y(_0882_));
NOR _2701_ (.A(_0860_),.B(_0882_),.Y(_0005_));
NOR _2702_ (.A(_1293_),.B(_1331_),.Y(_0883_));
NAND _2703_ (.A(\mem[10] [15]),.B(_1331_),.Y(_0884_));
NAND _2704_ (.A(_1333_),.B(_0884_),.Y(_0885_));
NOR _2705_ (.A(_0883_),.B(_0885_),.Y(_0886_));
NOR _2706_ (.A(_1308_),.B(_1331_),.Y(_0887_));
NAND _2707_ (.A(\mem[11] [15]),.B(_1331_),.Y(_0888_));
NAND _2708_ (.A(read_addr[0]),.B(_0888_),.Y(_0889_));
NOR _2709_ (.A(_0887_),.B(_0889_),.Y(_0890_));
NOR _2710_ (.A(_0886_),.B(_0890_),.Y(_0891_));
NOR _2711_ (.A(_1330_),.B(_0891_),.Y(_0892_));
NOR _2712_ (.A(_1331_),.B(\mem[7] [15]),.Y(_0893_));
NOR _2713_ (.A(read_addr[2]),.B(\mem[3] [15]),.Y(_0894_));
NOR _2714_ (.A(_0893_),.B(_0894_),.Y(_0895_));
NOR _2715_ (.A(_1333_),.B(_0895_),.Y(_0896_));
NOR _2716_ (.A(_1331_),.B(\mem[6] [15]),.Y(_0897_));
NOR _2717_ (.A(read_addr[2]),.B(\mem[2] [15]),.Y(_0898_));
NOR _2718_ (.A(_0897_),.B(_0898_),.Y(_0899_));
NOR _2719_ (.A(read_addr[0]),.B(_0899_),.Y(_0900_));
NOR _2720_ (.A(_0896_),.B(_0900_),.Y(_0901_));
NOR _2721_ (.A(read_addr[3]),.B(_0901_),.Y(_0902_));
NOR _2722_ (.A(_0892_),.B(_0902_),.Y(_0903_));
NOR _2723_ (.A(_1332_),.B(_0903_),.Y(_0904_));
NOR _2724_ (.A(read_addr[2]),.B(_1345_),.Y(_0905_));
NAND _2725_ (.A(\mem[12] [15]),.B(read_addr[2]),.Y(_0906_));
NAND _2726_ (.A(_1333_),.B(_0906_),.Y(_0907_));
NOR _2727_ (.A(_0905_),.B(_0907_),.Y(_0908_));
NOR _2728_ (.A(read_addr[2]),.B(_1346_),.Y(_0909_));
NAND _2729_ (.A(\mem[13] [15]),.B(read_addr[2]),.Y(_0910_));
NAND _2730_ (.A(read_addr[0]),.B(_0910_),.Y(_0911_));
NOR _2731_ (.A(_0909_),.B(_0911_),.Y(_0912_));
NOR _2732_ (.A(_0908_),.B(_0912_),.Y(_0913_));
NOR _2733_ (.A(_1330_),.B(_0913_),.Y(_0914_));
NOR _2734_ (.A(read_addr[2]),.B(\mem[1] [15]),.Y(_0915_));
NOR _2735_ (.A(_1331_),.B(\mem[5] [15]),.Y(_0916_));
NOR _2736_ (.A(_0915_),.B(_0916_),.Y(_0917_));
NOR _2737_ (.A(_1333_),.B(_0917_),.Y(_0918_));
NOR _2738_ (.A(read_addr[2]),.B(\mem[0] [15]),.Y(_0919_));
NOR _2739_ (.A(_1331_),.B(\mem[4] [15]),.Y(_0920_));
NOR _2740_ (.A(_0919_),.B(_0920_),.Y(_0921_));
NOR _2741_ (.A(read_addr[0]),.B(_0921_),.Y(_0922_));
NOR _2742_ (.A(_0918_),.B(_0922_),.Y(_0923_));
NOR _2743_ (.A(read_addr[3]),.B(_0923_),.Y(_0924_));
NOR _2744_ (.A(_0914_),.B(_0924_),.Y(_0925_));
NOR _2745_ (.A(read_addr[1]),.B(_0925_),.Y(_0926_));
NOR _2746_ (.A(_0904_),.B(_0926_),.Y(_0006_));
NOR _2747_ (.A(_1351_),.B(_1439_),.Y(_0927_));
NAND _2748_ (.A(_1352_),.B(_1440_),.Y(_0928_));
NOR _2749_ (.A(_1438_),.B(_0928_),.Y(_0929_));
NAND _2750_ (.A(_1437_),.B(_0927_),.Y(_0930_));
NOR _2751_ (.A(_1310_),.B(_0930_),.Y(_0931_));
NAND _2752_ (.A(we),.B(_0929_),.Y(_0932_));
NOR _2753_ (.A(data[0]),.B(_0932_),.Y(_0933_));
NOR _2754_ (.A(\mem[0] [0]),.B(_0931_),.Y(_0934_));
NOR _2755_ (.A(_0933_),.B(_0934_),.Y(_0016_));
NOR _2756_ (.A(data[1]),.B(_0932_),.Y(_0935_));
NOR _2757_ (.A(\mem[0] [1]),.B(_0931_),.Y(_0936_));
NOR _2758_ (.A(_0935_),.B(_0936_),.Y(_0023_));
NOR _2759_ (.A(data[2]),.B(_0932_),.Y(_0937_));
NOR _2760_ (.A(\mem[0] [2]),.B(_0931_),.Y(_0938_));
NOR _2761_ (.A(_0937_),.B(_0938_),.Y(_0024_));
NOR _2762_ (.A(data[3]),.B(_0932_),.Y(_0939_));
NOR _2763_ (.A(\mem[0] [3]),.B(_0931_),.Y(_0940_));
NOR _2764_ (.A(_0939_),.B(_0940_),.Y(_0025_));
NOR _2765_ (.A(data[4]),.B(_0932_),.Y(_0941_));
NOR _2766_ (.A(\mem[0] [4]),.B(_0931_),.Y(_0942_));
NOR _2767_ (.A(_0941_),.B(_0942_),.Y(_0026_));
NOR _2768_ (.A(data[5]),.B(_0932_),.Y(_0943_));
NOR _2769_ (.A(\mem[0] [5]),.B(_0931_),.Y(_0944_));
NOR _2770_ (.A(_0943_),.B(_0944_),.Y(_0027_));
NOR _2771_ (.A(data[6]),.B(_0932_),.Y(_0945_));
NOR _2772_ (.A(\mem[0] [6]),.B(_0931_),.Y(_0946_));
NOR _2773_ (.A(_0945_),.B(_0946_),.Y(_0028_));
NOR _2774_ (.A(data[7]),.B(_0932_),.Y(_0947_));
NOR _2775_ (.A(\mem[0] [7]),.B(_0931_),.Y(_0948_));
NOR _2776_ (.A(_0947_),.B(_0948_),.Y(_0029_));
NOR _2777_ (.A(data[8]),.B(_0932_),.Y(_0949_));
NOR _2778_ (.A(\mem[0] [8]),.B(_0931_),.Y(_0950_));
NOR _2779_ (.A(_0949_),.B(_0950_),.Y(_0030_));
NOR _2780_ (.A(data[9]),.B(_0932_),.Y(_0951_));
NOR _2781_ (.A(\mem[0] [9]),.B(_0931_),.Y(_0952_));
NOR _2782_ (.A(_0951_),.B(_0952_),.Y(_0031_));
NOR _2783_ (.A(data[10]),.B(_0932_),.Y(_0953_));
NOR _2784_ (.A(\mem[0] [10]),.B(_0931_),.Y(_0954_));
NOR _2785_ (.A(_0953_),.B(_0954_),.Y(_0017_));
NOR _2786_ (.A(data[11]),.B(_0932_),.Y(_0955_));
NOR _2787_ (.A(\mem[0] [11]),.B(_0931_),.Y(_0956_));
NOR _2788_ (.A(_0955_),.B(_0956_),.Y(_0018_));
NOR _2789_ (.A(data[12]),.B(_0932_),.Y(_0957_));
NOR _2790_ (.A(\mem[0] [12]),.B(_0931_),.Y(_0958_));
NOR _2791_ (.A(_0957_),.B(_0958_),.Y(_0019_));
NOR _2792_ (.A(data[13]),.B(_0932_),.Y(_0959_));
NOR _2793_ (.A(\mem[0] [13]),.B(_0931_),.Y(_0960_));
NOR _2794_ (.A(_0959_),.B(_0960_),.Y(_0020_));
NOR _2795_ (.A(data[14]),.B(_0932_),.Y(_0961_));
NOR _2796_ (.A(\mem[0] [14]),.B(_0931_),.Y(_0962_));
NOR _2797_ (.A(_0961_),.B(_0962_),.Y(_0021_));
NOR _2798_ (.A(data[15]),.B(_0932_),.Y(_0963_));
NOR _2799_ (.A(\mem[0] [15]),.B(_0931_),.Y(_0964_));
NOR _2800_ (.A(_0963_),.B(_0964_),.Y(_0022_));
NOR _2801_ (.A(_1478_),.B(_0928_),.Y(_0965_));
NAND _2802_ (.A(_1477_),.B(_0927_),.Y(_0966_));
NAND _2803_ (.A(_1402_),.B(_0965_),.Y(_0967_));
NAND _2804_ (.A(\mem[1] [0]),.B(_0966_),.Y(_0968_));
NAND _2805_ (.A(_0967_),.B(_0968_),.Y(_0128_));
NAND _2806_ (.A(_1405_),.B(_0965_),.Y(_0969_));
NAND _2807_ (.A(\mem[1] [1]),.B(_0966_),.Y(_0970_));
NAND _2808_ (.A(_0969_),.B(_0970_),.Y(_0135_));
NAND _2809_ (.A(_1408_),.B(_0965_),.Y(_0971_));
NAND _2810_ (.A(\mem[1] [2]),.B(_0966_),.Y(_0972_));
NAND _2811_ (.A(_0971_),.B(_0972_),.Y(_0136_));
NAND _2812_ (.A(_1357_),.B(_0965_),.Y(_0973_));
NAND _2813_ (.A(\mem[1] [3]),.B(_0966_),.Y(_0974_));
NAND _2814_ (.A(_0973_),.B(_0974_),.Y(_0137_));
NAND _2815_ (.A(_1361_),.B(_0965_),.Y(_0975_));
NAND _2816_ (.A(\mem[1] [4]),.B(_0966_),.Y(_0976_));
NAND _2817_ (.A(_0975_),.B(_0976_),.Y(_0138_));
NAND _2818_ (.A(_1364_),.B(_0965_),.Y(_0977_));
NAND _2819_ (.A(\mem[1] [5]),.B(_0966_),.Y(_0978_));
NAND _2820_ (.A(_0977_),.B(_0978_),.Y(_0139_));
NAND _2821_ (.A(_1367_),.B(_0965_),.Y(_0979_));
NAND _2822_ (.A(\mem[1] [6]),.B(_0966_),.Y(_0980_));
NAND _2823_ (.A(_0979_),.B(_0980_),.Y(_0140_));
NAND _2824_ (.A(_1370_),.B(_0965_),.Y(_0981_));
NAND _2825_ (.A(\mem[1] [7]),.B(_0966_),.Y(_0982_));
NAND _2826_ (.A(_0981_),.B(_0982_),.Y(_0141_));
NAND _2827_ (.A(_1372_),.B(_0965_),.Y(_0983_));
NAND _2828_ (.A(\mem[1] [8]),.B(_0966_),.Y(_0984_));
NAND _2829_ (.A(_0983_),.B(_0984_),.Y(_0142_));
NAND _2830_ (.A(_1375_),.B(_0965_),.Y(_0985_));
NAND _2831_ (.A(\mem[1] [9]),.B(_0966_),.Y(_0986_));
NAND _2832_ (.A(_0985_),.B(_0986_),.Y(_0143_));
NAND _2833_ (.A(_1379_),.B(_0965_),.Y(_0987_));
NAND _2834_ (.A(\mem[1] [10]),.B(_0966_),.Y(_0988_));
NAND _2835_ (.A(_0987_),.B(_0988_),.Y(_0129_));
NAND _2836_ (.A(_1382_),.B(_0965_),.Y(_0989_));
NAND _2837_ (.A(\mem[1] [11]),.B(_0966_),.Y(_0990_));
NAND _2838_ (.A(_0989_),.B(_0990_),.Y(_0130_));
NAND _2839_ (.A(_1385_),.B(_0965_),.Y(_0991_));
NAND _2840_ (.A(\mem[1] [12]),.B(_0966_),.Y(_0992_));
NAND _2841_ (.A(_0991_),.B(_0992_),.Y(_0131_));
NAND _2842_ (.A(_1388_),.B(_0965_),.Y(_0993_));
NAND _2843_ (.A(\mem[1] [13]),.B(_0966_),.Y(_0994_));
NAND _2844_ (.A(_0993_),.B(_0994_),.Y(_0132_));
NAND _2845_ (.A(_1391_),.B(_0965_),.Y(_0995_));
NAND _2846_ (.A(\mem[1] [14]),.B(_0966_),.Y(_0996_));
NAND _2847_ (.A(_0995_),.B(_0996_),.Y(_0133_));
NAND _2848_ (.A(_1393_),.B(_0965_),.Y(_0997_));
NAND _2849_ (.A(\mem[1] [15]),.B(_0966_),.Y(_0998_));
NAND _2850_ (.A(_0997_),.B(_0998_),.Y(_0134_));
NOR _2851_ (.A(_1350_),.B(_0928_),.Y(_0999_));
NAND _2852_ (.A(_1349_),.B(_0927_),.Y(_1000_));
NAND _2853_ (.A(_1402_),.B(_0999_),.Y(_1001_));
NAND _2854_ (.A(\mem[2] [0]),.B(_1000_),.Y(_1002_));
NAND _2855_ (.A(_1001_),.B(_1002_),.Y(_0144_));
NAND _2856_ (.A(_1405_),.B(_0999_),.Y(_1003_));
NAND _2857_ (.A(\mem[2] [1]),.B(_1000_),.Y(_1004_));
NAND _2858_ (.A(_1003_),.B(_1004_),.Y(_0151_));
NAND _2859_ (.A(_1408_),.B(_0999_),.Y(_1005_));
NAND _2860_ (.A(\mem[2] [2]),.B(_1000_),.Y(_1006_));
NAND _2861_ (.A(_1005_),.B(_1006_),.Y(_0152_));
NAND _2862_ (.A(_1357_),.B(_0999_),.Y(_1007_));
NAND _2863_ (.A(\mem[2] [3]),.B(_1000_),.Y(_1008_));
NAND _2864_ (.A(_1007_),.B(_1008_),.Y(_0153_));
NAND _2865_ (.A(_1361_),.B(_0999_),.Y(_1009_));
NAND _2866_ (.A(\mem[2] [4]),.B(_1000_),.Y(_1010_));
NAND _2867_ (.A(_1009_),.B(_1010_),.Y(_0154_));
NAND _2868_ (.A(_1364_),.B(_0999_),.Y(_1011_));
NAND _2869_ (.A(\mem[2] [5]),.B(_1000_),.Y(_1012_));
NAND _2870_ (.A(_1011_),.B(_1012_),.Y(_0155_));
NAND _2871_ (.A(_1367_),.B(_0999_),.Y(_1013_));
NAND _2872_ (.A(\mem[2] [6]),.B(_1000_),.Y(_1014_));
NAND _2873_ (.A(_1013_),.B(_1014_),.Y(_0156_));
NAND _2874_ (.A(_1370_),.B(_0999_),.Y(_1015_));
NAND _2875_ (.A(\mem[2] [7]),.B(_1000_),.Y(_1016_));
NAND _2876_ (.A(_1015_),.B(_1016_),.Y(_0157_));
NAND _2877_ (.A(_1372_),.B(_0999_),.Y(_1017_));
NAND _2878_ (.A(\mem[2] [8]),.B(_1000_),.Y(_1018_));
NAND _2879_ (.A(_1017_),.B(_1018_),.Y(_0158_));
NAND _2880_ (.A(_1375_),.B(_0999_),.Y(_1019_));
NAND _2881_ (.A(\mem[2] [9]),.B(_1000_),.Y(_1020_));
NAND _2882_ (.A(_1019_),.B(_1020_),.Y(_0159_));
NAND _2883_ (.A(_1379_),.B(_0999_),.Y(_1021_));
NAND _2884_ (.A(\mem[2] [10]),.B(_1000_),.Y(_1022_));
NAND _2885_ (.A(_1021_),.B(_1022_),.Y(_0145_));
NAND _2886_ (.A(_1382_),.B(_0999_),.Y(_1023_));
NAND _2887_ (.A(\mem[2] [11]),.B(_1000_),.Y(_1024_));
NAND _2888_ (.A(_1023_),.B(_1024_),.Y(_0146_));
NAND _2889_ (.A(_1385_),.B(_0999_),.Y(_1025_));
NAND _2890_ (.A(\mem[2] [12]),.B(_1000_),.Y(_1026_));
NAND _2891_ (.A(_1025_),.B(_1026_),.Y(_0147_));
NAND _2892_ (.A(_1388_),.B(_0999_),.Y(_1027_));
NAND _2893_ (.A(\mem[2] [13]),.B(_1000_),.Y(_1028_));
NAND _2894_ (.A(_1027_),.B(_1028_),.Y(_0148_));
NAND _2895_ (.A(_1391_),.B(_0999_),.Y(_1029_));
NAND _2896_ (.A(\mem[2] [14]),.B(_1000_),.Y(_1030_));
NAND _2897_ (.A(_1029_),.B(_1030_),.Y(_0149_));
NAND _2898_ (.A(_1393_),.B(_0999_),.Y(_1031_));
NAND _2899_ (.A(\mem[2] [15]),.B(_1000_),.Y(_1032_));
NAND _2900_ (.A(_1031_),.B(_1032_),.Y(_0150_));
NOR _2901_ (.A(_1399_),.B(_0928_),.Y(_1033_));
NAND _2902_ (.A(_1398_),.B(_0927_),.Y(_1034_));
NAND _2903_ (.A(_1402_),.B(_1033_),.Y(_1035_));
NAND _2904_ (.A(\mem[3] [0]),.B(_1034_),.Y(_1036_));
NAND _2905_ (.A(_1035_),.B(_1036_),.Y(_0160_));
NAND _2906_ (.A(_1405_),.B(_1033_),.Y(_1037_));
NAND _2907_ (.A(\mem[3] [1]),.B(_1034_),.Y(_1038_));
NAND _2908_ (.A(_1037_),.B(_1038_),.Y(_0167_));
NAND _2909_ (.A(_1408_),.B(_1033_),.Y(_1039_));
NAND _2910_ (.A(\mem[3] [2]),.B(_1034_),.Y(_1040_));
NAND _2911_ (.A(_1039_),.B(_1040_),.Y(_0168_));
NAND _2912_ (.A(_1357_),.B(_1033_),.Y(_1041_));
NAND _2913_ (.A(\mem[3] [3]),.B(_1034_),.Y(_1042_));
NAND _2914_ (.A(_1041_),.B(_1042_),.Y(_0169_));
NAND _2915_ (.A(_1361_),.B(_1033_),.Y(_1043_));
NAND _2916_ (.A(\mem[3] [4]),.B(_1034_),.Y(_1044_));
NAND _2917_ (.A(_1043_),.B(_1044_),.Y(_0170_));
NAND _2918_ (.A(_1364_),.B(_1033_),.Y(_1045_));
NAND _2919_ (.A(\mem[3] [5]),.B(_1034_),.Y(_1046_));
NAND _2920_ (.A(_1045_),.B(_1046_),.Y(_0171_));
NAND _2921_ (.A(_1367_),.B(_1033_),.Y(_1047_));
NAND _2922_ (.A(\mem[3] [6]),.B(_1034_),.Y(_1048_));
NAND _2923_ (.A(_1047_),.B(_1048_),.Y(_0172_));
NAND _2924_ (.A(_1370_),.B(_1033_),.Y(_1049_));
NAND _2925_ (.A(\mem[3] [7]),.B(_1034_),.Y(_1050_));
NAND _2926_ (.A(_1049_),.B(_1050_),.Y(_0173_));
NAND _2927_ (.A(_1372_),.B(_1033_),.Y(_1051_));
NAND _2928_ (.A(\mem[3] [8]),.B(_1034_),.Y(_1052_));
NAND _2929_ (.A(_1051_),.B(_1052_),.Y(_0174_));
NAND _2930_ (.A(_1375_),.B(_1033_),.Y(_1053_));
NAND _2931_ (.A(\mem[3] [9]),.B(_1034_),.Y(_1054_));
NAND _2932_ (.A(_1053_),.B(_1054_),.Y(_0175_));
NAND _2933_ (.A(_1379_),.B(_1033_),.Y(_1055_));
NAND _2934_ (.A(\mem[3] [10]),.B(_1034_),.Y(_1056_));
NAND _2935_ (.A(_1055_),.B(_1056_),.Y(_0161_));
NAND _2936_ (.A(_1382_),.B(_1033_),.Y(_1057_));
NAND _2937_ (.A(\mem[3] [11]),.B(_1034_),.Y(_1058_));
NAND _2938_ (.A(_1057_),.B(_1058_),.Y(_0162_));
NAND _2939_ (.A(_1385_),.B(_1033_),.Y(_1059_));
NAND _2940_ (.A(\mem[3] [12]),.B(_1034_),.Y(_1060_));
NAND _2941_ (.A(_1059_),.B(_1060_),.Y(_0163_));
NAND _2942_ (.A(_1388_),.B(_1033_),.Y(_1061_));
NAND _2943_ (.A(\mem[3] [13]),.B(_1034_),.Y(_1062_));
NAND _2944_ (.A(_1061_),.B(_1062_),.Y(_0164_));
NAND _2945_ (.A(_1391_),.B(_1033_),.Y(_1063_));
NAND _2946_ (.A(\mem[3] [14]),.B(_1034_),.Y(_1064_));
NAND _2947_ (.A(_1063_),.B(_1064_),.Y(_0165_));
NAND _2948_ (.A(_1393_),.B(_1033_),.Y(_1065_));
NAND _2949_ (.A(\mem[3] [15]),.B(_1034_),.Y(_1066_));
NAND _2950_ (.A(_1065_),.B(_1066_),.Y(_0166_));
NOR _2951_ (.A(write_addr[3]),.B(_1440_),.Y(_1067_));
NAND _2952_ (.A(_1313_),.B(_1439_),.Y(_1068_));
NOR _2953_ (.A(_1438_),.B(_1068_),.Y(_1069_));
NAND _2954_ (.A(_1437_),.B(_1067_),.Y(_1070_));
NAND _2955_ (.A(_1402_),.B(_1069_),.Y(_1071_));
NAND _2956_ (.A(\mem[4] [0]),.B(_1070_),.Y(_1072_));
NAND _2957_ (.A(_1071_),.B(_1072_),.Y(_0176_));
NAND _2958_ (.A(_1405_),.B(_1069_),.Y(_1073_));
NAND _2959_ (.A(\mem[4] [1]),.B(_1070_),.Y(_1074_));
NAND _2960_ (.A(_1073_),.B(_1074_),.Y(_0183_));
NAND _2961_ (.A(_1408_),.B(_1069_),.Y(_1075_));
NAND _2962_ (.A(\mem[4] [2]),.B(_1070_),.Y(_1076_));
NAND _2963_ (.A(_1075_),.B(_1076_),.Y(_0184_));
NAND _2964_ (.A(_1357_),.B(_1069_),.Y(_1077_));
NAND _2965_ (.A(\mem[4] [3]),.B(_1070_),.Y(_1078_));
NAND _2966_ (.A(_1077_),.B(_1078_),.Y(_0185_));
NAND _2967_ (.A(_1361_),.B(_1069_),.Y(_1079_));
NAND _2968_ (.A(\mem[4] [4]),.B(_1070_),.Y(_1080_));
NAND _2969_ (.A(_1079_),.B(_1080_),.Y(_0186_));
NAND _2970_ (.A(_1364_),.B(_1069_),.Y(_1081_));
NAND _2971_ (.A(\mem[4] [5]),.B(_1070_),.Y(_1082_));
NAND _2972_ (.A(_1081_),.B(_1082_),.Y(_0187_));
NAND _2973_ (.A(_1367_),.B(_1069_),.Y(_1083_));
NAND _2974_ (.A(\mem[4] [6]),.B(_1070_),.Y(_1084_));
NAND _2975_ (.A(_1083_),.B(_1084_),.Y(_0188_));
NAND _2976_ (.A(_1370_),.B(_1069_),.Y(_1085_));
NAND _2977_ (.A(\mem[4] [7]),.B(_1070_),.Y(_1086_));
NAND _2978_ (.A(_1085_),.B(_1086_),.Y(_0189_));
NAND _2979_ (.A(_1372_),.B(_1069_),.Y(_1087_));
NAND _2980_ (.A(\mem[4] [8]),.B(_1070_),.Y(_1088_));
NAND _2981_ (.A(_1087_),.B(_1088_),.Y(_0190_));
NAND _2982_ (.A(_1375_),.B(_1069_),.Y(_1089_));
NAND _2983_ (.A(\mem[4] [9]),.B(_1070_),.Y(_1090_));
NAND _2984_ (.A(_1089_),.B(_1090_),.Y(_0191_));
NAND _2985_ (.A(_1379_),.B(_1069_),.Y(_1091_));
NAND _2986_ (.A(\mem[4] [10]),.B(_1070_),.Y(_1092_));
NAND _2987_ (.A(_1091_),.B(_1092_),.Y(_0177_));
NAND _2988_ (.A(_1382_),.B(_1069_),.Y(_1093_));
NAND _2989_ (.A(\mem[4] [11]),.B(_1070_),.Y(_1094_));
NAND _2990_ (.A(_1093_),.B(_1094_),.Y(_0178_));
NAND _2991_ (.A(_1385_),.B(_1069_),.Y(_1095_));
NAND _2992_ (.A(\mem[4] [12]),.B(_1070_),.Y(_1096_));
NAND _2993_ (.A(_1095_),.B(_1096_),.Y(_0179_));
NAND _2994_ (.A(_1388_),.B(_1069_),.Y(_1097_));
NAND _2995_ (.A(\mem[4] [13]),.B(_1070_),.Y(_1098_));
NAND _2996_ (.A(_1097_),.B(_1098_),.Y(_0180_));
NAND _2997_ (.A(_1391_),.B(_1069_),.Y(_1099_));
NAND _2998_ (.A(\mem[4] [14]),.B(_1070_),.Y(_1100_));
NAND _2999_ (.A(_1099_),.B(_1100_),.Y(_0181_));
NAND _3000_ (.A(_1393_),.B(_1069_),.Y(_1101_));
NAND _3001_ (.A(\mem[4] [15]),.B(_1070_),.Y(_1102_));
NAND _3002_ (.A(_1101_),.B(_1102_),.Y(_0182_));
NOR _3003_ (.A(_1478_),.B(_1068_),.Y(_1103_));
NAND _3004_ (.A(_1477_),.B(_1067_),.Y(_1104_));
NAND _3005_ (.A(_1402_),.B(_1103_),.Y(_1105_));
NAND _3006_ (.A(\mem[5] [0]),.B(_1104_),.Y(_1106_));
NAND _3007_ (.A(_1105_),.B(_1106_),.Y(_0192_));
NAND _3008_ (.A(_1405_),.B(_1103_),.Y(_1107_));
NAND _3009_ (.A(\mem[5] [1]),.B(_1104_),.Y(_1108_));
NAND _3010_ (.A(_1107_),.B(_1108_),.Y(_0199_));
NAND _3011_ (.A(_1408_),.B(_1103_),.Y(_1109_));
NAND _3012_ (.A(\mem[5] [2]),.B(_1104_),.Y(_1110_));
NAND _3013_ (.A(_1109_),.B(_1110_),.Y(_0200_));
NAND _3014_ (.A(_1357_),.B(_1103_),.Y(_1111_));
NAND _3015_ (.A(\mem[5] [3]),.B(_1104_),.Y(_1112_));
NAND _3016_ (.A(_1111_),.B(_1112_),.Y(_0201_));
NAND _3017_ (.A(_1361_),.B(_1103_),.Y(_1113_));
NAND _3018_ (.A(\mem[5] [4]),.B(_1104_),.Y(_1114_));
NAND _3019_ (.A(_1113_),.B(_1114_),.Y(_0202_));
NAND _3020_ (.A(_1364_),.B(_1103_),.Y(_1115_));
NAND _3021_ (.A(\mem[5] [5]),.B(_1104_),.Y(_1116_));
NAND _3022_ (.A(_1115_),.B(_1116_),.Y(_0203_));
NAND _3023_ (.A(_1367_),.B(_1103_),.Y(_1117_));
NAND _3024_ (.A(\mem[5] [6]),.B(_1104_),.Y(_1118_));
NAND _3025_ (.A(_1117_),.B(_1118_),.Y(_0204_));
NAND _3026_ (.A(_1370_),.B(_1103_),.Y(_1119_));
NAND _3027_ (.A(\mem[5] [7]),.B(_1104_),.Y(_1120_));
NAND _3028_ (.A(_1119_),.B(_1120_),.Y(_0205_));
NAND _3029_ (.A(_1372_),.B(_1103_),.Y(_1121_));
NAND _3030_ (.A(\mem[5] [8]),.B(_1104_),.Y(_1122_));
NAND _3031_ (.A(_1121_),.B(_1122_),.Y(_0206_));
NAND _3032_ (.A(_1375_),.B(_1103_),.Y(_1123_));
NAND _3033_ (.A(\mem[5] [9]),.B(_1104_),.Y(_1124_));
NAND _3034_ (.A(_1123_),.B(_1124_),.Y(_0207_));
NAND _3035_ (.A(_1379_),.B(_1103_),.Y(_1125_));
NAND _3036_ (.A(\mem[5] [10]),.B(_1104_),.Y(_1126_));
NAND _3037_ (.A(_1125_),.B(_1126_),.Y(_0193_));
NAND _3038_ (.A(_1382_),.B(_1103_),.Y(_1127_));
NAND _3039_ (.A(\mem[5] [11]),.B(_1104_),.Y(_1128_));
NAND _3040_ (.A(_1127_),.B(_1128_),.Y(_0194_));
NAND _3041_ (.A(_1385_),.B(_1103_),.Y(_1129_));
NAND _3042_ (.A(\mem[5] [12]),.B(_1104_),.Y(_1130_));
NAND _3043_ (.A(_1129_),.B(_1130_),.Y(_0195_));
NAND _3044_ (.A(_1388_),.B(_1103_),.Y(_1131_));
NAND _3045_ (.A(\mem[5] [13]),.B(_1104_),.Y(_1132_));
NAND _3046_ (.A(_1131_),.B(_1132_),.Y(_0196_));
NAND _3047_ (.A(_1391_),.B(_1103_),.Y(_1133_));
NAND _3048_ (.A(\mem[5] [14]),.B(_1104_),.Y(_1134_));
NAND _3049_ (.A(_1133_),.B(_1134_),.Y(_0197_));
NAND _3050_ (.A(_1393_),.B(_1103_),.Y(_1135_));
NAND _3051_ (.A(\mem[5] [15]),.B(_1104_),.Y(_1136_));
NAND _3052_ (.A(_1135_),.B(_1136_),.Y(_0198_));
NOR _3053_ (.A(_1350_),.B(_1068_),.Y(_1137_));
NAND _3054_ (.A(_1349_),.B(_1067_),.Y(_1138_));
NAND _3055_ (.A(_1402_),.B(_1137_),.Y(_1139_));
NAND _3056_ (.A(\mem[6] [0]),.B(_1138_),.Y(_1140_));
NAND _3057_ (.A(_1139_),.B(_1140_),.Y(_0208_));
NAND _3058_ (.A(_1405_),.B(_1137_),.Y(_1141_));
NAND _3059_ (.A(\mem[6] [1]),.B(_1138_),.Y(_1142_));
NAND _3060_ (.A(_1141_),.B(_1142_),.Y(_0215_));
NAND _3061_ (.A(_1408_),.B(_1137_),.Y(_1143_));
NAND _3062_ (.A(\mem[6] [2]),.B(_1138_),.Y(_1144_));
NAND _3063_ (.A(_1143_),.B(_1144_),.Y(_0216_));
NAND _3064_ (.A(_1357_),.B(_1137_),.Y(_1145_));
NAND _3065_ (.A(\mem[6] [3]),.B(_1138_),.Y(_1146_));
NAND _3066_ (.A(_1145_),.B(_1146_),.Y(_0217_));
NAND _3067_ (.A(_1361_),.B(_1137_),.Y(_1147_));
NAND _3068_ (.A(\mem[6] [4]),.B(_1138_),.Y(_1148_));
NAND _3069_ (.A(_1147_),.B(_1148_),.Y(_0218_));
NAND _3070_ (.A(_1364_),.B(_1137_),.Y(_1149_));
NAND _3071_ (.A(\mem[6] [5]),.B(_1138_),.Y(_1150_));
NAND _3072_ (.A(_1149_),.B(_1150_),.Y(_0219_));
NAND _3073_ (.A(_1367_),.B(_1137_),.Y(_1151_));
NAND _3074_ (.A(\mem[6] [6]),.B(_1138_),.Y(_1152_));
NAND _3075_ (.A(_1151_),.B(_1152_),.Y(_0220_));
NAND _3076_ (.A(_1370_),.B(_1137_),.Y(_1153_));
NAND _3077_ (.A(\mem[6] [7]),.B(_1138_),.Y(_1154_));
NAND _3078_ (.A(_1153_),.B(_1154_),.Y(_0221_));
NAND _3079_ (.A(_1372_),.B(_1137_),.Y(_1155_));
NAND _3080_ (.A(\mem[6] [8]),.B(_1138_),.Y(_1156_));
NAND _3081_ (.A(_1155_),.B(_1156_),.Y(_0222_));
NAND _3082_ (.A(_1375_),.B(_1137_),.Y(_1157_));
NAND _3083_ (.A(\mem[6] [9]),.B(_1138_),.Y(_1158_));
NAND _3084_ (.A(_1157_),.B(_1158_),.Y(_0223_));
NAND _3085_ (.A(_1379_),.B(_1137_),.Y(_1159_));
NAND _3086_ (.A(\mem[6] [10]),.B(_1138_),.Y(_1160_));
NAND _3087_ (.A(_1159_),.B(_1160_),.Y(_0209_));
NAND _3088_ (.A(_1382_),.B(_1137_),.Y(_1161_));
NAND _3089_ (.A(\mem[6] [11]),.B(_1138_),.Y(_1162_));
NAND _3090_ (.A(_1161_),.B(_1162_),.Y(_0210_));
NAND _3091_ (.A(_1385_),.B(_1137_),.Y(_1163_));
NAND _3092_ (.A(\mem[6] [12]),.B(_1138_),.Y(_1164_));
NAND _3093_ (.A(_1163_),.B(_1164_),.Y(_0211_));
NAND _3094_ (.A(_1388_),.B(_1137_),.Y(_1165_));
NAND _3095_ (.A(\mem[6] [13]),.B(_1138_),.Y(_1166_));
NAND _3096_ (.A(_1165_),.B(_1166_),.Y(_0212_));
NAND _3097_ (.A(_1391_),.B(_1137_),.Y(_1167_));
NAND _3098_ (.A(\mem[6] [14]),.B(_1138_),.Y(_1168_));
NAND _3099_ (.A(_1167_),.B(_1168_),.Y(_0213_));
NAND _3100_ (.A(_1393_),.B(_1137_),.Y(_1169_));
NAND _3101_ (.A(\mem[6] [15]),.B(_1138_),.Y(_1170_));
NAND _3102_ (.A(_1169_),.B(_1170_),.Y(_0214_));
NOR _3103_ (.A(_1399_),.B(_1068_),.Y(_1171_));
NAND _3104_ (.A(_1398_),.B(_1067_),.Y(_1172_));
NAND _3105_ (.A(_1402_),.B(_1171_),.Y(_1173_));
NAND _3106_ (.A(\mem[7] [0]),.B(_1172_),.Y(_1174_));
NAND _3107_ (.A(_1173_),.B(_1174_),.Y(_0224_));
NAND _3108_ (.A(_1405_),.B(_1171_),.Y(_1175_));
NAND _3109_ (.A(\mem[7] [1]),.B(_1172_),.Y(_1176_));
NAND _3110_ (.A(_1175_),.B(_1176_),.Y(_0231_));
NAND _3111_ (.A(_1408_),.B(_1171_),.Y(_1177_));
NAND _3112_ (.A(\mem[7] [2]),.B(_1172_),.Y(_1178_));
NAND _3113_ (.A(_1177_),.B(_1178_),.Y(_0232_));
NAND _3114_ (.A(_1357_),.B(_1171_),.Y(_1179_));
NAND _3115_ (.A(\mem[7] [3]),.B(_1172_),.Y(_1180_));
NAND _3116_ (.A(_1179_),.B(_1180_),.Y(_0233_));
NAND _3117_ (.A(_1361_),.B(_1171_),.Y(_1181_));
NAND _3118_ (.A(\mem[7] [4]),.B(_1172_),.Y(_1182_));
NAND _3119_ (.A(_1181_),.B(_1182_),.Y(_0234_));
NAND _3120_ (.A(_1364_),.B(_1171_),.Y(_1183_));
NAND _3121_ (.A(\mem[7] [5]),.B(_1172_),.Y(_1184_));
NAND _3122_ (.A(_1183_),.B(_1184_),.Y(_0235_));
NAND _3123_ (.A(_1367_),.B(_1171_),.Y(_1185_));
NAND _3124_ (.A(\mem[7] [6]),.B(_1172_),.Y(_1186_));
NAND _3125_ (.A(_1185_),.B(_1186_),.Y(_0236_));
NAND _3126_ (.A(_1370_),.B(_1171_),.Y(_1187_));
NAND _3127_ (.A(\mem[7] [7]),.B(_1172_),.Y(_1188_));
NAND _3128_ (.A(_1187_),.B(_1188_),.Y(_0237_));
NAND _3129_ (.A(_1372_),.B(_1171_),.Y(_1189_));
NAND _3130_ (.A(\mem[7] [8]),.B(_1172_),.Y(_1190_));
NAND _3131_ (.A(_1189_),.B(_1190_),.Y(_0238_));
NAND _3132_ (.A(_1375_),.B(_1171_),.Y(_1191_));
NAND _3133_ (.A(\mem[7] [9]),.B(_1172_),.Y(_1192_));
NAND _3134_ (.A(_1191_),.B(_1192_),.Y(_0239_));
NAND _3135_ (.A(_1379_),.B(_1171_),.Y(_1193_));
NAND _3136_ (.A(\mem[7] [10]),.B(_1172_),.Y(_1194_));
NAND _3137_ (.A(_1193_),.B(_1194_),.Y(_0225_));
NAND _3138_ (.A(_1382_),.B(_1171_),.Y(_1195_));
NAND _3139_ (.A(\mem[7] [11]),.B(_1172_),.Y(_1196_));
NAND _3140_ (.A(_1195_),.B(_1196_),.Y(_0226_));
NAND _3141_ (.A(_1385_),.B(_1171_),.Y(_1197_));
NAND _3142_ (.A(\mem[7] [12]),.B(_1172_),.Y(_1198_));
NAND _3143_ (.A(_1197_),.B(_1198_),.Y(_0227_));
NAND _3144_ (.A(_1388_),.B(_1171_),.Y(_1199_));
NAND _3145_ (.A(\mem[7] [13]),.B(_1172_),.Y(_1200_));
NAND _3146_ (.A(_1199_),.B(_1200_),.Y(_0228_));
NAND _3147_ (.A(_1391_),.B(_1171_),.Y(_1201_));
NAND _3148_ (.A(\mem[7] [14]),.B(_1172_),.Y(_1202_));
NAND _3149_ (.A(_1201_),.B(_1202_),.Y(_0229_));
NAND _3150_ (.A(_1393_),.B(_1171_),.Y(_1203_));
NAND _3151_ (.A(\mem[7] [15]),.B(_1172_),.Y(_1204_));
NAND _3152_ (.A(_1203_),.B(_1204_),.Y(_0230_));
NOR _3153_ (.A(_1354_),.B(_1438_),.Y(_1205_));
NAND _3154_ (.A(_1353_),.B(_1437_),.Y(_1206_));
NAND _3155_ (.A(_1402_),.B(_1205_),.Y(_1207_));
NAND _3156_ (.A(\mem[8] [0]),.B(_1206_),.Y(_1208_));
NAND _3157_ (.A(_1207_),.B(_1208_),.Y(_0240_));
NAND _3158_ (.A(_1405_),.B(_1205_),.Y(_1209_));
NAND _3159_ (.A(\mem[8] [1]),.B(_1206_),.Y(_1210_));
NAND _3160_ (.A(_1209_),.B(_1210_),.Y(_0247_));
NAND _3161_ (.A(_1408_),.B(_1205_),.Y(_1211_));
NAND _3162_ (.A(\mem[8] [2]),.B(_1206_),.Y(_1212_));
NAND _3163_ (.A(_1211_),.B(_1212_),.Y(_0248_));
NAND _3164_ (.A(_1357_),.B(_1205_),.Y(_1213_));
NAND _3165_ (.A(\mem[8] [3]),.B(_1206_),.Y(_1214_));
NAND _3166_ (.A(_1213_),.B(_1214_),.Y(_0249_));
NAND _3167_ (.A(_1361_),.B(_1205_),.Y(_1215_));
NAND _3168_ (.A(\mem[8] [4]),.B(_1206_),.Y(_1216_));
NAND _3169_ (.A(_1215_),.B(_1216_),.Y(_0250_));
NAND _3170_ (.A(_1364_),.B(_1205_),.Y(_1217_));
NAND _3171_ (.A(\mem[8] [5]),.B(_1206_),.Y(_1218_));
NAND _3172_ (.A(_1217_),.B(_1218_),.Y(_0251_));
NAND _3173_ (.A(_1367_),.B(_1205_),.Y(_1219_));
NAND _3174_ (.A(\mem[8] [6]),.B(_1206_),.Y(_1220_));
NAND _3175_ (.A(_1219_),.B(_1220_),.Y(_0252_));
NAND _3176_ (.A(_1370_),.B(_1205_),.Y(_1221_));
NAND _3177_ (.A(\mem[8] [7]),.B(_1206_),.Y(_1222_));
NAND _3178_ (.A(_1221_),.B(_1222_),.Y(_0253_));
NAND _3179_ (.A(_1372_),.B(_1205_),.Y(_1223_));
NAND _3180_ (.A(\mem[8] [8]),.B(_1206_),.Y(_1224_));
NAND _3181_ (.A(_1223_),.B(_1224_),.Y(_0254_));
NAND _3182_ (.A(_1375_),.B(_1205_),.Y(_1225_));
NAND _3183_ (.A(\mem[8] [9]),.B(_1206_),.Y(_1226_));
NAND _3184_ (.A(_1225_),.B(_1226_),.Y(_0255_));
NAND _3185_ (.A(_1379_),.B(_1205_),.Y(_1227_));
NAND _3186_ (.A(\mem[8] [10]),.B(_1206_),.Y(_1228_));
NAND _3187_ (.A(_1227_),.B(_1228_),.Y(_0241_));
NAND _3188_ (.A(_1382_),.B(_1205_),.Y(_1229_));
NAND _3189_ (.A(\mem[8] [11]),.B(_1206_),.Y(_1230_));
NAND _3190_ (.A(_1229_),.B(_1230_),.Y(_0242_));
NAND _3191_ (.A(_1385_),.B(_1205_),.Y(_1231_));
NAND _3192_ (.A(\mem[8] [12]),.B(_1206_),.Y(_1232_));
NAND _3193_ (.A(_1231_),.B(_1232_),.Y(_0243_));
NAND _3194_ (.A(_1388_),.B(_1205_),.Y(_1233_));
NAND _3195_ (.A(\mem[8] [13]),.B(_1206_),.Y(_1234_));
NAND _3196_ (.A(_1233_),.B(_1234_),.Y(_0244_));
NAND _3197_ (.A(_1391_),.B(_1205_),.Y(_1235_));
NAND _3198_ (.A(\mem[8] [14]),.B(_1206_),.Y(_1236_));
NAND _3199_ (.A(_1235_),.B(_1236_),.Y(_0245_));
NAND _3200_ (.A(_1393_),.B(_1205_),.Y(_1237_));
NAND _3201_ (.A(\mem[8] [15]),.B(_1206_),.Y(_1238_));
NAND _3202_ (.A(_1237_),.B(_1238_),.Y(_0246_));
NOR _3203_ (.A(_1354_),.B(_1478_),.Y(_1239_));
NAND _3204_ (.A(_1353_),.B(_1477_),.Y(_1240_));
NAND _3205_ (.A(_1402_),.B(_1239_),.Y(_1241_));
NAND _3206_ (.A(\mem[9] [0]),.B(_1240_),.Y(_1242_));
NAND _3207_ (.A(_1241_),.B(_1242_),.Y(_0256_));
NAND _3208_ (.A(_1405_),.B(_1239_),.Y(_1243_));
NAND _3209_ (.A(\mem[9] [1]),.B(_1240_),.Y(_1244_));
NAND _3210_ (.A(_1243_),.B(_1244_),.Y(_0263_));
NAND _3211_ (.A(_1408_),.B(_1239_),.Y(_1245_));
NAND _3212_ (.A(\mem[9] [2]),.B(_1240_),.Y(_1246_));
NAND _3213_ (.A(_1245_),.B(_1246_),.Y(_0264_));
NAND _3214_ (.A(_1357_),.B(_1239_),.Y(_1247_));
NAND _3215_ (.A(\mem[9] [3]),.B(_1240_),.Y(_1248_));
NAND _3216_ (.A(_1247_),.B(_1248_),.Y(_0265_));
NAND _3217_ (.A(_1361_),.B(_1239_),.Y(_1249_));
NAND _3218_ (.A(\mem[9] [4]),.B(_1240_),.Y(_1250_));
NAND _3219_ (.A(_1249_),.B(_1250_),.Y(_0266_));
NAND _3220_ (.A(_1364_),.B(_1239_),.Y(_1251_));
NAND _3221_ (.A(\mem[9] [5]),.B(_1240_),.Y(_1252_));
NAND _3222_ (.A(_1251_),.B(_1252_),.Y(_0267_));
NAND _3223_ (.A(_1367_),.B(_1239_),.Y(_1253_));
NAND _3224_ (.A(\mem[9] [6]),.B(_1240_),.Y(_1254_));
NAND _3225_ (.A(_1253_),.B(_1254_),.Y(_0268_));
NAND _3226_ (.A(_1370_),.B(_1239_),.Y(_1255_));
NAND _3227_ (.A(\mem[9] [7]),.B(_1240_),.Y(_1256_));
NAND _3228_ (.A(_1255_),.B(_1256_),.Y(_0269_));
NAND _3229_ (.A(_1372_),.B(_1239_),.Y(_1257_));
NAND _3230_ (.A(\mem[9] [8]),.B(_1240_),.Y(_1258_));
NAND _3231_ (.A(_1257_),.B(_1258_),.Y(_0270_));
NAND _3232_ (.A(_1375_),.B(_1239_),.Y(_1259_));
NAND _3233_ (.A(\mem[9] [9]),.B(_1240_),.Y(_1260_));
NAND _3234_ (.A(_1259_),.B(_1260_),.Y(_0271_));
NAND _3235_ (.A(_1379_),.B(_1239_),.Y(_1261_));
NAND _3236_ (.A(\mem[9] [10]),.B(_1240_),.Y(_1262_));
NAND _3237_ (.A(_1261_),.B(_1262_),.Y(_0257_));
NAND _3238_ (.A(_1382_),.B(_1239_),.Y(_1263_));
NAND _3239_ (.A(\mem[9] [11]),.B(_1240_),.Y(_1264_));
NAND _3240_ (.A(_1263_),.B(_1264_),.Y(_0258_));
NAND _3241_ (.A(_1385_),.B(_1239_),.Y(_1265_));
NAND _3242_ (.A(\mem[9] [12]),.B(_1240_),.Y(_1266_));
NAND _3243_ (.A(_1265_),.B(_1266_),.Y(_0259_));
NAND _3244_ (.A(_1388_),.B(_1239_),.Y(_1267_));
NAND _3245_ (.A(\mem[9] [13]),.B(_1240_),.Y(_1268_));
NAND _3246_ (.A(_1267_),.B(_1268_),.Y(_0260_));
NAND _3247_ (.A(_1391_),.B(_1239_),.Y(_1269_));
NAND _3248_ (.A(\mem[9] [14]),.B(_1240_),.Y(_1270_));
NAND _3249_ (.A(_1269_),.B(_1270_),.Y(_0261_));
NAND _3250_ (.A(_1393_),.B(_1239_),.Y(_1271_));
NAND _3251_ (.A(\mem[9] [15]),.B(_1240_),.Y(_1272_));
NAND _3252_ (.A(_1271_),.B(_1272_),.Y(_0262_));
NAND _3253_ (.A(_1355_),.B(_1402_),.Y(_1273_));
NAND _3254_ (.A(\mem[10] [0]),.B(_1356_),.Y(_1274_));
NAND _3255_ (.A(_1273_),.B(_1274_),.Y(_0032_));
NAND _3256_ (.A(\mem[10] [1]),.B(_1356_),.Y(_1275_));
NAND _3257_ (.A(_1355_),.B(_1405_),.Y(_1276_));
NAND _3258_ (.A(_1275_),.B(_1276_),.Y(_0039_));
NAND _3259_ (.A(\mem[10] [2]),.B(_1356_),.Y(_1277_));
NAND _3260_ (.A(_1355_),.B(_1408_),.Y(_1278_));
NAND _3261_ (.A(_1277_),.B(_1278_),.Y(_0040_));
DFF _3262_ (.C(write_clk),.D(_0016_),.Q(\mem[0] [0]));
DFF _3263_ (.C(write_clk),.D(_0023_),.Q(\mem[0] [1]));
DFF _3264_ (.C(write_clk),.D(_0024_),.Q(\mem[0] [2]));
DFF _3265_ (.C(write_clk),.D(_0025_),.Q(\mem[0] [3]));
DFF _3266_ (.C(write_clk),.D(_0026_),.Q(\mem[0] [4]));
DFF _3267_ (.C(write_clk),.D(_0027_),.Q(\mem[0] [5]));
DFF _3268_ (.C(write_clk),.D(_0028_),.Q(\mem[0] [6]));
DFF _3269_ (.C(write_clk),.D(_0029_),.Q(\mem[0] [7]));
DFF _3270_ (.C(write_clk),.D(_0030_),.Q(\mem[0] [8]));
DFF _3271_ (.C(write_clk),.D(_0031_),.Q(\mem[0] [9]));
DFF _3272_ (.C(write_clk),.D(_0017_),.Q(\mem[0] [10]));
DFF _3273_ (.C(write_clk),.D(_0018_),.Q(\mem[0] [11]));
DFF _3274_ (.C(write_clk),.D(_0019_),.Q(\mem[0] [12]));
DFF _3275_ (.C(write_clk),.D(_0020_),.Q(\mem[0] [13]));
DFF _3276_ (.C(write_clk),.D(_0021_),.Q(\mem[0] [14]));
DFF _3277_ (.C(write_clk),.D(_0022_),.Q(\mem[0] [15]));
DFF _3278_ (.C(write_clk),.D(_0144_),.Q(\mem[2] [0]));
DFF _3279_ (.C(write_clk),.D(_0151_),.Q(\mem[2] [1]));
DFF _3280_ (.C(write_clk),.D(_0152_),.Q(\mem[2] [2]));
DFF _3281_ (.C(write_clk),.D(_0153_),.Q(\mem[2] [3]));
DFF _3282_ (.C(write_clk),.D(_0154_),.Q(\mem[2] [4]));
DFF _3283_ (.C(write_clk),.D(_0155_),.Q(\mem[2] [5]));
DFF _3284_ (.C(write_clk),.D(_0156_),.Q(\mem[2] [6]));
DFF _3285_ (.C(write_clk),.D(_0157_),.Q(\mem[2] [7]));
DFF _3286_ (.C(write_clk),.D(_0158_),.Q(\mem[2] [8]));
DFF _3287_ (.C(write_clk),.D(_0159_),.Q(\mem[2] [9]));
DFF _3288_ (.C(write_clk),.D(_0145_),.Q(\mem[2] [10]));
DFF _3289_ (.C(write_clk),.D(_0146_),.Q(\mem[2] [11]));
DFF _3290_ (.C(write_clk),.D(_0147_),.Q(\mem[2] [12]));
DFF _3291_ (.C(write_clk),.D(_0148_),.Q(\mem[2] [13]));
DFF _3292_ (.C(write_clk),.D(_0149_),.Q(\mem[2] [14]));
DFF _3293_ (.C(write_clk),.D(_0150_),.Q(\mem[2] [15]));
DFF _3294_ (.C(write_clk),.D(_0176_),.Q(\mem[4] [0]));
DFF _3295_ (.C(write_clk),.D(_0183_),.Q(\mem[4] [1]));
DFF _3296_ (.C(write_clk),.D(_0184_),.Q(\mem[4] [2]));
DFF _3297_ (.C(write_clk),.D(_0185_),.Q(\mem[4] [3]));
DFF _3298_ (.C(write_clk),.D(_0186_),.Q(\mem[4] [4]));
DFF _3299_ (.C(write_clk),.D(_0187_),.Q(\mem[4] [5]));
DFF _3300_ (.C(write_clk),.D(_0188_),.Q(\mem[4] [6]));
DFF _3301_ (.C(write_clk),.D(_0189_),.Q(\mem[4] [7]));
DFF _3302_ (.C(write_clk),.D(_0190_),.Q(\mem[4] [8]));
DFF _3303_ (.C(write_clk),.D(_0191_),.Q(\mem[4] [9]));
DFF _3304_ (.C(write_clk),.D(_0177_),.Q(\mem[4] [10]));
DFF _3305_ (.C(write_clk),.D(_0178_),.Q(\mem[4] [11]));
DFF _3306_ (.C(write_clk),.D(_0179_),.Q(\mem[4] [12]));
DFF _3307_ (.C(write_clk),.D(_0180_),.Q(\mem[4] [13]));
DFF _3308_ (.C(write_clk),.D(_0181_),.Q(\mem[4] [14]));
DFF _3309_ (.C(write_clk),.D(_0182_),.Q(\mem[4] [15]));
DFF _3310_ (.C(write_clk),.D(_0160_),.Q(\mem[3] [0]));
DFF _3311_ (.C(write_clk),.D(_0167_),.Q(\mem[3] [1]));
DFF _3312_ (.C(write_clk),.D(_0168_),.Q(\mem[3] [2]));
DFF _3313_ (.C(write_clk),.D(_0169_),.Q(\mem[3] [3]));
DFF _3314_ (.C(write_clk),.D(_0170_),.Q(\mem[3] [4]));
DFF _3315_ (.C(write_clk),.D(_0171_),.Q(\mem[3] [5]));
DFF _3316_ (.C(write_clk),.D(_0172_),.Q(\mem[3] [6]));
DFF _3317_ (.C(write_clk),.D(_0173_),.Q(\mem[3] [7]));
DFF _3318_ (.C(write_clk),.D(_0174_),.Q(\mem[3] [8]));
DFF _3319_ (.C(write_clk),.D(_0175_),.Q(\mem[3] [9]));
DFF _3320_ (.C(write_clk),.D(_0161_),.Q(\mem[3] [10]));
DFF _3321_ (.C(write_clk),.D(_0162_),.Q(\mem[3] [11]));
DFF _3322_ (.C(write_clk),.D(_0163_),.Q(\mem[3] [12]));
DFF _3323_ (.C(write_clk),.D(_0164_),.Q(\mem[3] [13]));
DFF _3324_ (.C(write_clk),.D(_0165_),.Q(\mem[3] [14]));
DFF _3325_ (.C(write_clk),.D(_0166_),.Q(\mem[3] [15]));
DFF _3326_ (.C(write_clk),.D(_0128_),.Q(\mem[1] [0]));
DFF _3327_ (.C(write_clk),.D(_0135_),.Q(\mem[1] [1]));
DFF _3328_ (.C(write_clk),.D(_0136_),.Q(\mem[1] [2]));
DFF _3329_ (.C(write_clk),.D(_0137_),.Q(\mem[1] [3]));
DFF _3330_ (.C(write_clk),.D(_0138_),.Q(\mem[1] [4]));
DFF _3331_ (.C(write_clk),.D(_0139_),.Q(\mem[1] [5]));
DFF _3332_ (.C(write_clk),.D(_0140_),.Q(\mem[1] [6]));
DFF _3333_ (.C(write_clk),.D(_0141_),.Q(\mem[1] [7]));
DFF _3334_ (.C(write_clk),.D(_0142_),.Q(\mem[1] [8]));
DFF _3335_ (.C(write_clk),.D(_0143_),.Q(\mem[1] [9]));
DFF _3336_ (.C(write_clk),.D(_0129_),.Q(\mem[1] [10]));
DFF _3337_ (.C(write_clk),.D(_0130_),.Q(\mem[1] [11]));
DFF _3338_ (.C(write_clk),.D(_0131_),.Q(\mem[1] [12]));
DFF _3339_ (.C(write_clk),.D(_0132_),.Q(\mem[1] [13]));
DFF _3340_ (.C(write_clk),.D(_0133_),.Q(\mem[1] [14]));
DFF _3341_ (.C(write_clk),.D(_0134_),.Q(\mem[1] [15]));
DFF _3342_ (.C(write_clk),.D(_0192_),.Q(\mem[5] [0]));
DFF _3343_ (.C(write_clk),.D(_0199_),.Q(\mem[5] [1]));
DFF _3344_ (.C(write_clk),.D(_0200_),.Q(\mem[5] [2]));
DFF _3345_ (.C(write_clk),.D(_0201_),.Q(\mem[5] [3]));
DFF _3346_ (.C(write_clk),.D(_0202_),.Q(\mem[5] [4]));
DFF _3347_ (.C(write_clk),.D(_0203_),.Q(\mem[5] [5]));
DFF _3348_ (.C(write_clk),.D(_0204_),.Q(\mem[5] [6]));
DFF _3349_ (.C(write_clk),.D(_0205_),.Q(\mem[5] [7]));
DFF _3350_ (.C(write_clk),.D(_0206_),.Q(\mem[5] [8]));
DFF _3351_ (.C(write_clk),.D(_0207_),.Q(\mem[5] [9]));
DFF _3352_ (.C(write_clk),.D(_0193_),.Q(\mem[5] [10]));
DFF _3353_ (.C(write_clk),.D(_0194_),.Q(\mem[5] [11]));
DFF _3354_ (.C(write_clk),.D(_0195_),.Q(\mem[5] [12]));
DFF _3355_ (.C(write_clk),.D(_0196_),.Q(\mem[5] [13]));
DFF _3356_ (.C(write_clk),.D(_0197_),.Q(\mem[5] [14]));
DFF _3357_ (.C(write_clk),.D(_0198_),.Q(\mem[5] [15]));
DFF _3358_ (.C(write_clk),.D(_0208_),.Q(\mem[6] [0]));
DFF _3359_ (.C(write_clk),.D(_0215_),.Q(\mem[6] [1]));
DFF _3360_ (.C(write_clk),.D(_0216_),.Q(\mem[6] [2]));
DFF _3361_ (.C(write_clk),.D(_0217_),.Q(\mem[6] [3]));
DFF _3362_ (.C(write_clk),.D(_0218_),.Q(\mem[6] [4]));
DFF _3363_ (.C(write_clk),.D(_0219_),.Q(\mem[6] [5]));
DFF _3364_ (.C(write_clk),.D(_0220_),.Q(\mem[6] [6]));
DFF _3365_ (.C(write_clk),.D(_0221_),.Q(\mem[6] [7]));
DFF _3366_ (.C(write_clk),.D(_0222_),.Q(\mem[6] [8]));
DFF _3367_ (.C(write_clk),.D(_0223_),.Q(\mem[6] [9]));
DFF _3368_ (.C(write_clk),.D(_0209_),.Q(\mem[6] [10]));
DFF _3369_ (.C(write_clk),.D(_0210_),.Q(\mem[6] [11]));
DFF _3370_ (.C(write_clk),.D(_0211_),.Q(\mem[6] [12]));
DFF _3371_ (.C(write_clk),.D(_0212_),.Q(\mem[6] [13]));
DFF _3372_ (.C(write_clk),.D(_0213_),.Q(\mem[6] [14]));
DFF _3373_ (.C(write_clk),.D(_0214_),.Q(\mem[6] [15]));
DFF _3374_ (.C(write_clk),.D(_0224_),.Q(\mem[7] [0]));
DFF _3375_ (.C(write_clk),.D(_0231_),.Q(\mem[7] [1]));
DFF _3376_ (.C(write_clk),.D(_0232_),.Q(\mem[7] [2]));
DFF _3377_ (.C(write_clk),.D(_0233_),.Q(\mem[7] [3]));
DFF _3378_ (.C(write_clk),.D(_0234_),.Q(\mem[7] [4]));
DFF _3379_ (.C(write_clk),.D(_0235_),.Q(\mem[7] [5]));
DFF _3380_ (.C(write_clk),.D(_0236_),.Q(\mem[7] [6]));
DFF _3381_ (.C(write_clk),.D(_0237_),.Q(\mem[7] [7]));
DFF _3382_ (.C(write_clk),.D(_0238_),.Q(\mem[7] [8]));
DFF _3383_ (.C(write_clk),.D(_0239_),.Q(\mem[7] [9]));
DFF _3384_ (.C(write_clk),.D(_0225_),.Q(\mem[7] [10]));
DFF _3385_ (.C(write_clk),.D(_0226_),.Q(\mem[7] [11]));
DFF _3386_ (.C(write_clk),.D(_0227_),.Q(\mem[7] [12]));
DFF _3387_ (.C(write_clk),.D(_0228_),.Q(\mem[7] [13]));
DFF _3388_ (.C(write_clk),.D(_0229_),.Q(\mem[7] [14]));
DFF _3389_ (.C(write_clk),.D(_0230_),.Q(\mem[7] [15]));
DFF _3390_ (.C(write_clk),.D(_0240_),.Q(\mem[8] [0]));
DFF _3391_ (.C(write_clk),.D(_0247_),.Q(\mem[8] [1]));
DFF _3392_ (.C(write_clk),.D(_0248_),.Q(\mem[8] [2]));
DFF _3393_ (.C(write_clk),.D(_0249_),.Q(\mem[8] [3]));
DFF _3394_ (.C(write_clk),.D(_0250_),.Q(\mem[8] [4]));
DFF _3395_ (.C(write_clk),.D(_0251_),.Q(\mem[8] [5]));
DFF _3396_ (.C(write_clk),.D(_0252_),.Q(\mem[8] [6]));
DFF _3397_ (.C(write_clk),.D(_0253_),.Q(\mem[8] [7]));
DFF _3398_ (.C(write_clk),.D(_0254_),.Q(\mem[8] [8]));
DFF _3399_ (.C(write_clk),.D(_0255_),.Q(\mem[8] [9]));
DFF _3400_ (.C(write_clk),.D(_0241_),.Q(\mem[8] [10]));
DFF _3401_ (.C(write_clk),.D(_0242_),.Q(\mem[8] [11]));
DFF _3402_ (.C(write_clk),.D(_0243_),.Q(\mem[8] [12]));
DFF _3403_ (.C(write_clk),.D(_0244_),.Q(\mem[8] [13]));
DFF _3404_ (.C(write_clk),.D(_0245_),.Q(\mem[8] [14]));
DFF _3405_ (.C(write_clk),.D(_0246_),.Q(\mem[8] [15]));
DFF _3406_ (.C(write_clk),.D(_0256_),.Q(\mem[9] [0]));
DFF _3407_ (.C(write_clk),.D(_0263_),.Q(\mem[9] [1]));
DFF _3408_ (.C(write_clk),.D(_0264_),.Q(\mem[9] [2]));
DFF _3409_ (.C(write_clk),.D(_0265_),.Q(\mem[9] [3]));
DFF _3410_ (.C(write_clk),.D(_0266_),.Q(\mem[9] [4]));
DFF _3411_ (.C(write_clk),.D(_0267_),.Q(\mem[9] [5]));
DFF _3412_ (.C(write_clk),.D(_0268_),.Q(\mem[9] [6]));
DFF _3413_ (.C(write_clk),.D(_0269_),.Q(\mem[9] [7]));
DFF _3414_ (.C(write_clk),.D(_0270_),.Q(\mem[9] [8]));
DFF _3415_ (.C(write_clk),.D(_0271_),.Q(\mem[9] [9]));
DFF _3416_ (.C(write_clk),.D(_0257_),.Q(\mem[9] [10]));
DFF _3417_ (.C(write_clk),.D(_0258_),.Q(\mem[9] [11]));
DFF _3418_ (.C(write_clk),.D(_0259_),.Q(\mem[9] [12]));
DFF _3419_ (.C(write_clk),.D(_0260_),.Q(\mem[9] [13]));
DFF _3420_ (.C(write_clk),.D(_0261_),.Q(\mem[9] [14]));
DFF _3421_ (.C(write_clk),.D(_0262_),.Q(\mem[9] [15]));
DFF _3422_ (.C(write_clk),.D(_0032_),.Q(\mem[10] [0]));
DFF _3423_ (.C(write_clk),.D(_0039_),.Q(\mem[10] [1]));
DFF _3424_ (.C(write_clk),.D(_0040_),.Q(\mem[10] [2]));
DFF _3425_ (.C(write_clk),.D(_0041_),.Q(\mem[10] [3]));
DFF _3426_ (.C(write_clk),.D(_0042_),.Q(\mem[10] [4]));
DFF _3427_ (.C(write_clk),.D(_0043_),.Q(\mem[10] [5]));
DFF _3428_ (.C(write_clk),.D(_0044_),.Q(\mem[10] [6]));
DFF _3429_ (.C(write_clk),.D(_0045_),.Q(\mem[10] [7]));
DFF _3430_ (.C(write_clk),.D(_0046_),.Q(\mem[10] [8]));
DFF _3431_ (.C(write_clk),.D(_0047_),.Q(\mem[10] [9]));
DFF _3432_ (.C(write_clk),.D(_0033_),.Q(\mem[10] [10]));
DFF _3433_ (.C(write_clk),.D(_0034_),.Q(\mem[10] [11]));
DFF _3434_ (.C(write_clk),.D(_0035_),.Q(\mem[10] [12]));
DFF _3435_ (.C(write_clk),.D(_0036_),.Q(\mem[10] [13]));
DFF _3436_ (.C(write_clk),.D(_0037_),.Q(\mem[10] [14]));
DFF _3437_ (.C(write_clk),.D(_0038_),.Q(\mem[10] [15]));
DFF _3438_ (.C(write_clk),.D(_0048_),.Q(\mem[11] [0]));
DFF _3439_ (.C(write_clk),.D(_0055_),.Q(\mem[11] [1]));
DFF _3440_ (.C(write_clk),.D(_0056_),.Q(\mem[11] [2]));
DFF _3441_ (.C(write_clk),.D(_0057_),.Q(\mem[11] [3]));
DFF _3442_ (.C(write_clk),.D(_0058_),.Q(\mem[11] [4]));
DFF _3443_ (.C(write_clk),.D(_0059_),.Q(\mem[11] [5]));
DFF _3444_ (.C(write_clk),.D(_0060_),.Q(\mem[11] [6]));
DFF _3445_ (.C(write_clk),.D(_0061_),.Q(\mem[11] [7]));
DFF _3446_ (.C(write_clk),.D(_0062_),.Q(\mem[11] [8]));
DFF _3447_ (.C(write_clk),.D(_0063_),.Q(\mem[11] [9]));
DFF _3448_ (.C(write_clk),.D(_0049_),.Q(\mem[11] [10]));
DFF _3449_ (.C(write_clk),.D(_0050_),.Q(\mem[11] [11]));
DFF _3450_ (.C(write_clk),.D(_0051_),.Q(\mem[11] [12]));
DFF _3451_ (.C(write_clk),.D(_0052_),.Q(\mem[11] [13]));
DFF _3452_ (.C(write_clk),.D(_0053_),.Q(\mem[11] [14]));
DFF _3453_ (.C(write_clk),.D(_0054_),.Q(\mem[11] [15]));
DFF _3454_ (.C(write_clk),.D(_0064_),.Q(\mem[12] [0]));
DFF _3455_ (.C(write_clk),.D(_0071_),.Q(\mem[12] [1]));
DFF _3456_ (.C(write_clk),.D(_0072_),.Q(\mem[12] [2]));
DFF _3457_ (.C(write_clk),.D(_0073_),.Q(\mem[12] [3]));
DFF _3458_ (.C(write_clk),.D(_0074_),.Q(\mem[12] [4]));
DFF _3459_ (.C(write_clk),.D(_0075_),.Q(\mem[12] [5]));
DFF _3460_ (.C(write_clk),.D(_0076_),.Q(\mem[12] [6]));
DFF _3461_ (.C(write_clk),.D(_0077_),.Q(\mem[12] [7]));
DFF _3462_ (.C(write_clk),.D(_0078_),.Q(\mem[12] [8]));
DFF _3463_ (.C(write_clk),.D(_0079_),.Q(\mem[12] [9]));
DFF _3464_ (.C(write_clk),.D(_0065_),.Q(\mem[12] [10]));
DFF _3465_ (.C(write_clk),.D(_0066_),.Q(\mem[12] [11]));
DFF _3466_ (.C(write_clk),.D(_0067_),.Q(\mem[12] [12]));
DFF _3467_ (.C(write_clk),.D(_0068_),.Q(\mem[12] [13]));
DFF _3468_ (.C(write_clk),.D(_0069_),.Q(\mem[12] [14]));
DFF _3469_ (.C(write_clk),.D(_0070_),.Q(\mem[12] [15]));
DFF _3470_ (.C(write_clk),.D(_0080_),.Q(\mem[13] [0]));
DFF _3471_ (.C(write_clk),.D(_0087_),.Q(\mem[13] [1]));
DFF _3472_ (.C(write_clk),.D(_0088_),.Q(\mem[13] [2]));
DFF _3473_ (.C(write_clk),.D(_0089_),.Q(\mem[13] [3]));
DFF _3474_ (.C(write_clk),.D(_0090_),.Q(\mem[13] [4]));
DFF _3475_ (.C(write_clk),.D(_0091_),.Q(\mem[13] [5]));
DFF _3476_ (.C(write_clk),.D(_0092_),.Q(\mem[13] [6]));
DFF _3477_ (.C(write_clk),.D(_0093_),.Q(\mem[13] [7]));
DFF _3478_ (.C(write_clk),.D(_0094_),.Q(\mem[13] [8]));
DFF _3479_ (.C(write_clk),.D(_0095_),.Q(\mem[13] [9]));
DFF _3480_ (.C(write_clk),.D(_0081_),.Q(\mem[13] [10]));
DFF _3481_ (.C(write_clk),.D(_0082_),.Q(\mem[13] [11]));
DFF _3482_ (.C(write_clk),.D(_0083_),.Q(\mem[13] [12]));
DFF _3483_ (.C(write_clk),.D(_0084_),.Q(\mem[13] [13]));
DFF _3484_ (.C(write_clk),.D(_0085_),.Q(\mem[13] [14]));
DFF _3485_ (.C(write_clk),.D(_0086_),.Q(\mem[13] [15]));
DFF _3486_ (.C(write_clk),.D(_0096_),.Q(\mem[14] [0]));
DFF _3487_ (.C(write_clk),.D(_0103_),.Q(\mem[14] [1]));
DFF _3488_ (.C(write_clk),.D(_0104_),.Q(\mem[14] [2]));
DFF _3489_ (.C(write_clk),.D(_0105_),.Q(\mem[14] [3]));
DFF _3490_ (.C(write_clk),.D(_0106_),.Q(\mem[14] [4]));
DFF _3491_ (.C(write_clk),.D(_0107_),.Q(\mem[14] [5]));
DFF _3492_ (.C(write_clk),.D(_0108_),.Q(\mem[14] [6]));
DFF _3493_ (.C(write_clk),.D(_0109_),.Q(\mem[14] [7]));
DFF _3494_ (.C(write_clk),.D(_0110_),.Q(\mem[14] [8]));
DFF _3495_ (.C(write_clk),.D(_0111_),.Q(\mem[14] [9]));
DFF _3496_ (.C(write_clk),.D(_0097_),.Q(\mem[14] [10]));
DFF _3497_ (.C(write_clk),.D(_0098_),.Q(\mem[14] [11]));
DFF _3498_ (.C(write_clk),.D(_0099_),.Q(\mem[14] [12]));
DFF _3499_ (.C(write_clk),.D(_0100_),.Q(\mem[14] [13]));
DFF _3500_ (.C(write_clk),.D(_0101_),.Q(\mem[14] [14]));
DFF _3501_ (.C(write_clk),.D(_0102_),.Q(\mem[14] [15]));
DFF _3502_ (.C(write_clk),.D(_0112_),.Q(\mem[15] [0]));
DFF _3503_ (.C(write_clk),.D(_0119_),.Q(\mem[15] [1]));
DFF _3504_ (.C(write_clk),.D(_0120_),.Q(\mem[15] [2]));
DFF _3505_ (.C(write_clk),.D(_0121_),.Q(\mem[15] [3]));
DFF _3506_ (.C(write_clk),.D(_0122_),.Q(\mem[15] [4]));
DFF _3507_ (.C(write_clk),.D(_0123_),.Q(\mem[15] [5]));
DFF _3508_ (.C(write_clk),.D(_0124_),.Q(\mem[15] [6]));
DFF _3509_ (.C(write_clk),.D(_0125_),.Q(\mem[15] [7]));
DFF _3510_ (.C(write_clk),.D(_0126_),.Q(\mem[15] [8]));
DFF _3511_ (.C(write_clk),.D(_0127_),.Q(\mem[15] [9]));
DFF _3512_ (.C(write_clk),.D(_0113_),.Q(\mem[15] [10]));
DFF _3513_ (.C(write_clk),.D(_0114_),.Q(\mem[15] [11]));
DFF _3514_ (.C(write_clk),.D(_0115_),.Q(\mem[15] [12]));
DFF _3515_ (.C(write_clk),.D(_0116_),.Q(\mem[15] [13]));
DFF _3516_ (.C(write_clk),.D(_0117_),.Q(\mem[15] [14]));
DFF _3517_ (.C(write_clk),.D(_0118_),.Q(\mem[15] [15]));
DFF _3518_ (.C(read_clk),.D(_0000_),.Q(q[0]));
DFF _3519_ (.C(read_clk),.D(_0007_),.Q(q[1]));
DFF _3520_ (.C(read_clk),.D(_0008_),.Q(q[2]));
DFF _3521_ (.C(read_clk),.D(_0009_),.Q(q[3]));
DFF _3522_ (.C(read_clk),.D(_0010_),.Q(q[4]));
DFF _3523_ (.C(read_clk),.D(_0011_),.Q(q[5]));
DFF _3524_ (.C(read_clk),.D(_0012_),.Q(q[6]));
DFF _3525_ (.C(read_clk),.D(_0013_),.Q(q[7]));
DFF _3526_ (.C(read_clk),.D(_0014_),.Q(q[8]));
DFF _3527_ (.C(read_clk),.D(_0015_),.Q(q[9]));
DFF _3528_ (.C(read_clk),.D(_0001_),.Q(q[10]));
DFF _3529_ (.C(read_clk),.D(_0002_),.Q(q[11]));
DFF _3530_ (.C(read_clk),.D(_0003_),.Q(q[12]));
DFF _3531_ (.C(read_clk),.D(_0004_),.Q(q[13]));
DFF _3532_ (.C(read_clk),.D(_0005_),.Q(q[14]));
DFF _3533_ (.C(read_clk),.D(_0006_),.Q(q[15]));
endmodule